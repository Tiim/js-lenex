<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Schwimmclub Fricktal" version="11.70661">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Frick" name="Fricktal-Cup" course="SCM" deadline="2021-09-10" entrystartdate="2021-07-12" entrytype="INVITATION" hostclub="Schwimmclub Fricktal" hostclub.url="http://www.scfricktal.ch" number="14" organizer="SCFTAL" organizer.url="http://www.scfricktal.ch/" reservecount="2" result.url="https://live.swimrankings.net/29421/" startmethod="1" timing="AUTOMATIC" type="SUI.IM" withdrawuntil="2021-09-10" state="AG" nation="SUI">
      <AGEDATE value="2021-01-01" type="YEAR" />
      <POOL name="Hallenbad Rain, 5070 Frick" lanemin="1" lanemax="4" />
      <FACILITY city="Frick" name="Hallenbad Rain, 5070 Frick" nation="SUI" state="AG" street="Juraweg 13" zip="5070" />
      <POINTTABLE pointtableid="3014" name="FINA Point Scoring" version="2021" />
      <CONTACT city="5070" email="meldungen@scfricktal.ch" name="Schwimmclub Fricktal" street="Hallenbad Rain" street2="Juraweg 13" zip="Frick" />
      <FEES>
        <FEE currency="CHF" type="LATEENTRY.INDIVIDUAL" value="500" />
        <FEE currency="CHF" type="LATEENTRY.RELAY" value="1000" />
      </FEES>
      <SESSIONS>
        <SESSION date="2021-09-18" daytime="08:30" endtime="12:30" name="Vormittag" number="1" officialmeeting="08:00" teamleadermeeting="07:45" warmupfrom="07:30" warmupuntil="08:15">
          <EVENTS>
            <EVENT eventid="1053" daytime="08:30" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1056" agemax="9" agemin="-1" name="9 Jahre und jünger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12342" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1057" agemax="10" agemin="10" name="10 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14229" />
                    <RANKING order="2" place="-1" resultid="14279" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1058" agemax="11" agemin="11" name="11 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13477" />
                    <RANKING order="2" place="2" resultid="13481" />
                    <RANKING order="3" place="3" resultid="13470" />
                    <RANKING order="4" place="4" resultid="13082" />
                    <RANKING order="5" place="5" resultid="13191" />
                    <RANKING order="6" place="6" resultid="14342" />
                    <RANKING order="7" place="7" resultid="14243" />
                    <RANKING order="8" place="-1" resultid="13106" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1055" agemax="12" agemin="12" name="12 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13536" />
                    <RANKING order="2" place="2" resultid="13451" />
                    <RANKING order="3" place="3" resultid="14521" />
                    <RANKING order="4" place="4" resultid="14533" />
                    <RANKING order="5" place="5" resultid="13492" />
                    <RANKING order="6" place="6" resultid="14556" />
                    <RANKING order="7" place="7" resultid="13666" />
                    <RANKING order="8" place="8" resultid="14275" />
                    <RANKING order="9" place="9" resultid="14635" />
                    <RANKING order="10" place="10" resultid="12355" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12846" daytime="08:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12847" daytime="08:31" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12848" daytime="08:33" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="12849" daytime="08:34" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="12850" daytime="08:35" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="12851" daytime="08:37" number="6" order="6" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="*" timestandardlistid="5603">
                  <FEE currency="CHF" value="1000" />
                </TIMESTANDARDREF>
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1060" daytime="08:38" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1061" agemax="9" agemin="-1" name="9 Jahre und jünger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14304" />
                    <RANKING order="2" place="2" resultid="14208" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1062" agemax="10" agemin="10" name="10 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12385" />
                    <RANKING order="2" place="-1" resultid="12445" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1063" agemax="11" agemin="11" name="11 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12441" />
                    <RANKING order="2" place="2" resultid="12380" />
                    <RANKING order="3" place="3" resultid="14263" />
                    <RANKING order="4" place="-1" resultid="14320" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1064" agemax="12" agemin="12" name="12 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13194" />
                    <RANKING order="2" place="2" resultid="12450" />
                    <RANKING order="3" place="3" resultid="13213" />
                    <RANKING order="4" place="4" resultid="14548" />
                    <RANKING order="5" place="5" resultid="12351" />
                    <RANKING order="6" place="6" resultid="14117" />
                    <RANKING order="7" place="-1" resultid="14611" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12852" daytime="08:38" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12853" daytime="08:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12854" daytime="08:41" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="12855" daytime="08:42" number="4" order="4" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="*" timestandardlistid="5601">
                  <FEE currency="CHF" value="1000" />
                </TIMESTANDARDREF>
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1065" daytime="08:44" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1066" agemax="11" agemin="11" name="11 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14575" />
                    <RANKING order="2" place="2" resultid="14591" />
                    <RANKING order="3" place="3" resultid="13482" />
                    <RANKING order="4" place="4" resultid="13698" />
                    <RANKING order="5" place="5" resultid="13083" />
                    <RANKING order="6" place="6" resultid="13241" />
                    <RANKING order="7" place="7" resultid="13192" />
                    <RANKING order="8" place="8" resultid="14583" />
                    <RANKING order="9" place="9" resultid="14126" />
                    <RANKING order="10" place="10" resultid="14188" />
                    <RANKING order="11" place="11" resultid="14200" />
                    <RANKING order="12" place="12" resultid="14240" />
                    <RANKING order="13" place="-1" resultid="13447" />
                    <RANKING order="14" place="-1" resultid="13425" />
                    <RANKING order="15" place="-1" resultid="13222" />
                    <RANKING order="16" place="-1" resultid="13107" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1067" agemax="12" agemin="12" name="12 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14537" />
                    <RANKING order="2" place="2" resultid="13459" />
                    <RANKING order="3" place="3" resultid="13526" />
                    <RANKING order="4" place="4" resultid="14276" />
                    <RANKING order="5" place="5" resultid="14615" />
                    <RANKING order="6" place="6" resultid="14164" />
                    <RANKING order="7" place="7" resultid="14131" />
                    <RANKING order="8" place="8" resultid="14639" />
                    <RANKING order="9" place="9" resultid="13691" />
                    <RANKING order="10" place="10" resultid="13735" />
                    <RANKING order="11" place="11" resultid="12401" />
                    <RANKING order="12" place="12" resultid="12356" />
                    <RANKING order="13" place="13" resultid="12364" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12856" daytime="08:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12857" daytime="08:47" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12858" daytime="08:49" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="12859" daytime="08:52" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="12860" daytime="08:54" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="12861" daytime="08:56" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="12862" daytime="08:58" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="12863" daytime="09:00" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1070" daytime="09:03" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1071" agemax="11" agemin="11" name="11 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14571" />
                    <RANKING order="2" place="2" resultid="13455" />
                    <RANKING order="3" place="3" resultid="12442" />
                    <RANKING order="4" place="4" resultid="12347" />
                    <RANKING order="5" place="5" resultid="12381" />
                    <RANKING order="6" place="6" resultid="13154" />
                    <RANKING order="7" place="7" resultid="13443" />
                    <RANKING order="8" place="8" resultid="13233" />
                    <RANKING order="9" place="9" resultid="14323" />
                    <RANKING order="10" place="10" resultid="12405" />
                    <RANKING order="11" place="11" resultid="13437" />
                    <RANKING order="12" place="-1" resultid="14309" />
                    <RANKING order="13" place="-1" resultid="12413" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1072" agemax="12" agemin="12" name="12 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13195" />
                    <RANKING order="2" place="2" resultid="13709" />
                    <RANKING order="3" place="3" resultid="13226" />
                    <RANKING order="4" place="4" resultid="13214" />
                    <RANKING order="5" place="5" resultid="13653" />
                    <RANKING order="6" place="6" resultid="14118" />
                    <RANKING order="7" place="-1" resultid="14529" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12864" daytime="09:03" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12865" daytime="09:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12866" daytime="09:08" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="12867" daytime="09:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="12868" daytime="09:12" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1073" daytime="09:15" gender="F" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1074" agemax="9" agemin="-1" name="9 Jahre und jünger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12360" />
                    <RANKING order="2" place="2" resultid="14204" />
                    <RANKING order="3" place="3" resultid="14254" />
                    <RANKING order="4" place="4" resultid="13132" />
                    <RANKING order="5" place="5" resultid="13677" />
                    <RANKING order="6" place="6" resultid="13732" />
                    <RANKING order="7" place="7" resultid="12343" />
                    <RANKING order="8" place="8" resultid="12389" />
                    <RANKING order="9" place="9" resultid="14292" />
                    <RANKING order="10" place="10" resultid="14329" />
                    <RANKING order="11" place="11" resultid="14222" />
                    <RANKING order="12" place="-1" resultid="14284" />
                    <RANKING order="13" place="-1" resultid="14338" />
                    <RANKING order="14" place="-1" resultid="14245" />
                    <RANKING order="15" place="-1" resultid="14213" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1075" agemax="10" agemin="10" name="10 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13649" />
                    <RANKING order="2" place="2" resultid="14139" />
                    <RANKING order="3" place="3" resultid="13102" />
                    <RANKING order="4" place="4" resultid="13661" />
                    <RANKING order="5" place="5" resultid="14236" />
                    <RANKING order="6" place="6" resultid="14184" />
                    <RANKING order="7" place="7" resultid="13180" />
                    <RANKING order="8" place="8" resultid="13502" />
                    <RANKING order="9" place="9" resultid="14226" />
                    <RANKING order="10" place="10" resultid="13127" />
                    <RANKING order="11" place="11" resultid="13097" />
                    <RANKING order="12" place="12" resultid="13673" />
                    <RANKING order="13" place="13" resultid="13062" />
                    <RANKING order="14" place="-1" resultid="14272" />
                    <RANKING order="15" place="-1" resultid="13058" />
                    <RANKING order="16" place="-1" resultid="14280" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12870" daytime="09:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12871" daytime="09:17" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12872" daytime="09:19" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="12873" daytime="09:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="12874" daytime="09:22" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="12875" daytime="09:23" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="12876" daytime="09:24" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="12877" daytime="09:26" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1076" daytime="09:28" gender="M" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1077" agemax="9" agemin="-1" name="9 Jahre und jünger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13237" />
                    <RANKING order="2" place="2" resultid="14305" />
                    <RANKING order="3" place="3" resultid="14209" />
                    <RANKING order="4" place="4" resultid="13078" />
                    <RANKING order="5" place="5" resultid="14325" />
                    <RANKING order="6" place="6" resultid="14122" />
                    <RANKING order="7" place="7" resultid="12454" />
                    <RANKING order="8" place="8" resultid="13631" />
                    <RANKING order="9" place="9" resultid="13218" />
                    <RANKING order="10" place="-1" resultid="14150" />
                    <RANKING order="11" place="-1" resultid="14268" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1078" agemax="10" agemin="10" name="10 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12446" />
                    <RANKING order="2" place="2" resultid="12437" />
                    <RANKING order="3" place="3" resultid="13123" />
                    <RANKING order="4" place="4" resultid="13093" />
                    <RANKING order="5" place="5" resultid="14143" />
                    <RANKING order="6" place="6" resultid="13634" />
                    <RANKING order="7" place="-1" resultid="14296" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12878" daytime="09:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12879" daytime="09:29" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12880" daytime="09:31" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="12881" daytime="09:33" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="12882" daytime="09:34" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1084" daytime="09:36" gender="F" number="7" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1085" agemax="10" agemin="10" name="10 Jahre" />
                <AGEGROUP agegroupid="1087" agemax="11" agemin="11" name="11 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14343" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1086" agemax="12" agemin="12" name="12 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13493" />
                    <RANKING order="2" place="2" resultid="13452" />
                    <RANKING order="3" place="3" resultid="13537" />
                    <RANKING order="4" place="4" resultid="14147" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12883" daytime="09:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="14112" daytime="09:40" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="*" timestandardlistid="5603">
                  <FEE currency="CHF" value="1000" />
                </TIMESTANDARDREF>
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1088" daytime="09:43" gender="M" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1089" agemax="10" agemin="10" name="10 Jahre" />
                <AGEGROUP agegroupid="1090" agemax="11" agemin="11" name="11 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14264" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1091" agemax="12" agemin="12" name="12 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12451" />
                    <RANKING order="2" place="2" resultid="13216" />
                    <RANKING order="3" place="3" resultid="12352" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12884" daytime="09:43" number="1" order="1" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="*" timestandardlistid="5601">
                  <FEE currency="CHF" value="1000" />
                </TIMESTANDARDREF>
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1092" daytime="09:48" gender="F" number="9" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1093" agemax="9" agemin="-1" name="9 Jahre und jünger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12344" />
                    <RANKING order="2" place="2" resultid="14255" />
                    <RANKING order="3" place="3" resultid="14339" />
                    <RANKING order="4" place="4" resultid="14205" />
                    <RANKING order="5" place="5" resultid="12361" />
                    <RANKING order="6" place="6" resultid="12390" />
                    <RANKING order="7" place="7" resultid="14293" />
                    <RANKING order="8" place="8" resultid="13133" />
                    <RANKING order="9" place="9" resultid="14330" />
                    <RANKING order="10" place="10" resultid="14285" />
                    <RANKING order="11" place="11" resultid="14223" />
                    <RANKING order="12" place="-1" resultid="14246" />
                    <RANKING order="13" place="-1" resultid="14214" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1094" agemax="10" agemin="10" name="10 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13650" />
                    <RANKING order="2" place="2" resultid="13662" />
                    <RANKING order="3" place="3" resultid="14140" />
                    <RANKING order="4" place="4" resultid="14237" />
                    <RANKING order="5" place="5" resultid="13503" />
                    <RANKING order="6" place="6" resultid="13128" />
                    <RANKING order="7" place="7" resultid="14227" />
                    <RANKING order="8" place="8" resultid="13098" />
                    <RANKING order="9" place="9" resultid="13103" />
                    <RANKING order="10" place="10" resultid="14185" />
                    <RANKING order="11" place="11" resultid="13674" />
                    <RANKING order="12" place="-1" resultid="13063" />
                    <RANKING order="13" place="-1" resultid="13181" />
                    <RANKING order="14" place="-1" resultid="14273" />
                    <RANKING order="15" place="-1" resultid="13059" />
                    <RANKING order="16" place="-1" resultid="14281" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12885" daytime="09:48" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12886" daytime="09:49" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12887" daytime="09:51" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="12888" daytime="09:53" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="12889" daytime="09:54" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="12890" daytime="09:56" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="12891" daytime="09:57" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="14113" daytime="09:59" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1096" daytime="10:01" gender="M" number="10" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1097" agemax="9" agemin="-1" name="9 Jahre und jünger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13238" />
                    <RANKING order="2" place="2" resultid="14306" />
                    <RANKING order="3" place="3" resultid="14123" />
                    <RANKING order="4" place="4" resultid="13219" />
                    <RANKING order="5" place="5" resultid="14210" />
                    <RANKING order="6" place="6" resultid="13079" />
                    <RANKING order="7" place="7" resultid="14326" />
                    <RANKING order="8" place="-1" resultid="14151" />
                    <RANKING order="9" place="-1" resultid="12455" />
                    <RANKING order="10" place="-1" resultid="14269" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1098" agemax="10" agemin="10" name="10 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12438" />
                    <RANKING order="2" place="2" resultid="13094" />
                    <RANKING order="3" place="3" resultid="12447" />
                    <RANKING order="4" place="4" resultid="12386" />
                    <RANKING order="5" place="5" resultid="13124" />
                    <RANKING order="6" place="6" resultid="14144" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12892" daytime="10:01" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12893" daytime="10:03" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12894" daytime="10:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="12895" daytime="10:06" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1099" daytime="10:08" gender="F" number="11" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1102" agemax="11" agemin="11" name="11 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14576" />
                    <RANKING order="2" place="2" resultid="13471" />
                    <RANKING order="3" place="3" resultid="14584" />
                    <RANKING order="4" place="4" resultid="13448" />
                    <RANKING order="5" place="5" resultid="13478" />
                    <RANKING order="6" place="6" resultid="14592" />
                    <RANKING order="7" place="7" resultid="13699" />
                    <RANKING order="8" place="8" resultid="13084" />
                    <RANKING order="9" place="9" resultid="13243" />
                    <RANKING order="10" place="10" resultid="13223" />
                    <RANKING order="11" place="11" resultid="14127" />
                    <RANKING order="12" place="12" resultid="13189" />
                    <RANKING order="13" place="13" resultid="14201" />
                    <RANKING order="14" place="14" resultid="14241" />
                    <RANKING order="15" place="-1" resultid="13108" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1101" agemax="12" agemin="12" name="12 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14522" />
                    <RANKING order="2" place="2" resultid="13665" />
                    <RANKING order="3" place="3" resultid="14534" />
                    <RANKING order="4" place="4" resultid="13460" />
                    <RANKING order="5" place="5" resultid="14165" />
                    <RANKING order="6" place="6" resultid="14636" />
                    <RANKING order="7" place="7" resultid="14640" />
                    <RANKING order="8" place="8" resultid="14557" />
                    <RANKING order="9" place="9" resultid="14564" />
                    <RANKING order="10" place="10" resultid="14616" />
                    <RANKING order="11" place="11" resultid="13736" />
                    <RANKING order="12" place="12" resultid="14130" />
                    <RANKING order="13" place="13" resultid="13692" />
                    <RANKING order="14" place="14" resultid="12365" />
                    <RANKING order="15" place="15" resultid="12402" />
                    <RANKING order="16" place="-1" resultid="13527" />
                    <RANKING order="17" place="-1" resultid="12357" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12897" daytime="10:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12898" daytime="10:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12899" daytime="10:13" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="12900" daytime="10:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="12901" daytime="10:18" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="12902" daytime="10:20" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="12903" daytime="10:22" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="12904" daytime="10:24" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1103" daytime="10:27" gender="M" number="12" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1104" agemax="11" agemin="11" name="11 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14572" />
                    <RANKING order="2" place="2" resultid="12348" />
                    <RANKING order="3" place="3" resultid="13456" />
                    <RANKING order="4" place="4" resultid="12382" />
                    <RANKING order="5" place="5" resultid="13234" />
                    <RANKING order="6" place="6" resultid="14321" />
                    <RANKING order="7" place="7" resultid="14265" />
                    <RANKING order="8" place="8" resultid="13546" />
                    <RANKING order="9" place="9" resultid="13155" />
                    <RANKING order="10" place="-1" resultid="12406" />
                    <RANKING order="11" place="-1" resultid="12414" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1105" agemax="12" agemin="12" name="12 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14549" />
                    <RANKING order="2" place="2" resultid="13196" />
                    <RANKING order="3" place="3" resultid="13710" />
                    <RANKING order="4" place="4" resultid="14530" />
                    <RANKING order="5" place="5" resultid="13654" />
                    <RANKING order="6" place="6" resultid="14612" />
                    <RANKING order="7" place="7" resultid="14119" />
                    <RANKING order="8" place="-1" resultid="13533" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12906" daytime="10:27" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12907" daytime="10:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12908" daytime="10:32" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="12909" daytime="10:35" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="12910" daytime="10:37" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1106" daytime="10:40" gender="F" number="13" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1107" agemax="9" agemin="-1" name="9 Jahre und jünger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12345" />
                    <RANKING order="2" place="2" resultid="12362" />
                    <RANKING order="3" place="3" resultid="13134" />
                    <RANKING order="4" place="4" resultid="14206" />
                    <RANKING order="5" place="5" resultid="12391" />
                    <RANKING order="6" place="6" resultid="13678" />
                    <RANKING order="7" place="7" resultid="14256" />
                    <RANKING order="8" place="8" resultid="13733" />
                    <RANKING order="9" place="9" resultid="14294" />
                    <RANKING order="10" place="10" resultid="14340" />
                    <RANKING order="11" place="11" resultid="14286" />
                    <RANKING order="12" place="12" resultid="14331" />
                    <RANKING order="13" place="13" resultid="14247" />
                    <RANKING order="14" place="14" resultid="14224" />
                    <RANKING order="15" place="15" resultid="14215" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1108" agemax="10" agemin="10" name="10 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13651" />
                    <RANKING order="2" place="2" resultid="13104" />
                    <RANKING order="3" place="3" resultid="14141" />
                    <RANKING order="4" place="4" resultid="13182" />
                    <RANKING order="5" place="5" resultid="13504" />
                    <RANKING order="6" place="6" resultid="14228" />
                    <RANKING order="7" place="7" resultid="14186" />
                    <RANKING order="8" place="8" resultid="13099" />
                    <RANKING order="9" place="9" resultid="13129" />
                    <RANKING order="10" place="10" resultid="13663" />
                    <RANKING order="11" place="11" resultid="14238" />
                    <RANKING order="12" place="12" resultid="13675" />
                    <RANKING order="13" place="13" resultid="13064" />
                    <RANKING order="14" place="-1" resultid="13060" />
                    <RANKING order="15" place="-1" resultid="14282" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12911" daytime="10:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12912" daytime="10:42" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12913" daytime="10:43" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="12914" daytime="10:45" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="12915" daytime="10:46" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="12916" daytime="10:47" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="12917" daytime="10:49" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="12918" daytime="10:50" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1109" daytime="10:52" gender="M" number="14" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1110" agemax="9" agemin="-1" name="9 Jahre und jünger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14211" />
                    <RANKING order="2" place="2" resultid="13239" />
                    <RANKING order="3" place="3" resultid="14307" />
                    <RANKING order="4" place="4" resultid="13080" />
                    <RANKING order="5" place="5" resultid="14327" />
                    <RANKING order="6" place="6" resultid="14152" />
                    <RANKING order="7" place="7" resultid="14124" />
                    <RANKING order="8" place="8" resultid="13220" />
                    <RANKING order="9" place="9" resultid="12456" />
                    <RANKING order="10" place="10" resultid="13632" />
                    <RANKING order="11" place="11" resultid="14270" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1111" agemax="10" agemin="10" name="10 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12439" />
                    <RANKING order="2" place="2" resultid="12448" />
                    <RANKING order="3" place="3" resultid="13125" />
                    <RANKING order="4" place="4" resultid="13095" />
                    <RANKING order="5" place="5" resultid="14145" />
                    <RANKING order="6" place="6" resultid="13635" />
                    <RANKING order="7" place="7" resultid="14297" />
                    <RANKING order="8" place="-1" resultid="12387" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12919" daytime="10:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12920" daytime="10:53" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12921" daytime="10:55" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="12922" daytime="10:56" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="12923" daytime="10:57" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1112" daytime="10:59" gender="F" number="15" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1115" agemax="11" agemin="11" name="11 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14577" />
                    <RANKING order="2" place="2" resultid="13472" />
                    <RANKING order="3" place="3" resultid="13700" />
                    <RANKING order="4" place="4" resultid="14593" />
                    <RANKING order="5" place="5" resultid="13479" />
                    <RANKING order="6" place="6" resultid="13190" />
                    <RANKING order="7" place="7" resultid="13483" />
                    <RANKING order="8" place="8" resultid="13085" />
                    <RANKING order="9" place="9" resultid="13449" />
                    <RANKING order="10" place="10" resultid="14585" />
                    <RANKING order="11" place="11" resultid="13242" />
                    <RANKING order="12" place="12" resultid="13426" />
                    <RANKING order="13" place="13" resultid="14344" />
                    <RANKING order="14" place="14" resultid="14189" />
                    <RANKING order="15" place="15" resultid="14128" />
                    <RANKING order="16" place="16" resultid="13224" />
                    <RANKING order="17" place="17" resultid="14202" />
                    <RANKING order="18" place="18" resultid="14242" />
                    <RANKING order="19" place="-1" resultid="13109" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1114" agemax="12" agemin="12" name="12 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14538" />
                    <RANKING order="2" place="2" resultid="14523" />
                    <RANKING order="3" place="3" resultid="13494" />
                    <RANKING order="4" place="4" resultid="13453" />
                    <RANKING order="5" place="5" resultid="14535" />
                    <RANKING order="6" place="6" resultid="13538" />
                    <RANKING order="7" place="7" resultid="13461" />
                    <RANKING order="8" place="8" resultid="13667" />
                    <RANKING order="9" place="9" resultid="13528" />
                    <RANKING order="10" place="10" resultid="14277" />
                    <RANKING order="11" place="11" resultid="14637" />
                    <RANKING order="12" place="12" resultid="14148" />
                    <RANKING order="13" place="13" resultid="14558" />
                    <RANKING order="14" place="14" resultid="14617" />
                    <RANKING order="15" place="15" resultid="14565" />
                    <RANKING order="16" place="16" resultid="12403" />
                    <RANKING order="17" place="17" resultid="13737" />
                    <RANKING order="18" place="18" resultid="14166" />
                    <RANKING order="19" place="19" resultid="13693" />
                    <RANKING order="20" place="20" resultid="14641" />
                    <RANKING order="21" place="21" resultid="12358" />
                    <RANKING order="22" place="22" resultid="14132" />
                    <RANKING order="23" place="23" resultid="12366" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12925" daytime="10:59" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12926" daytime="11:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12927" daytime="11:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="12928" daytime="11:06" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="12929" daytime="11:08" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="12930" daytime="11:10" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="12931" daytime="11:12" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="12932" daytime="11:14" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="12933" daytime="11:16" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="12934" daytime="11:18" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="12935" daytime="11:20" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1116" daytime="11:22" gender="M" number="16" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1117" agemax="11" agemin="11" name="11 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14573" />
                    <RANKING order="2" place="2" resultid="12349" />
                    <RANKING order="3" place="3" resultid="13457" />
                    <RANKING order="4" place="4" resultid="12443" />
                    <RANKING order="5" place="5" resultid="12383" />
                    <RANKING order="6" place="6" resultid="13235" />
                    <RANKING order="7" place="7" resultid="13156" />
                    <RANKING order="8" place="8" resultid="12407" />
                    <RANKING order="9" place="9" resultid="14266" />
                    <RANKING order="10" place="10" resultid="13444" />
                    <RANKING order="11" place="11" resultid="14322" />
                    <RANKING order="12" place="12" resultid="13438" />
                    <RANKING order="13" place="13" resultid="13547" />
                    <RANKING order="14" place="-1" resultid="12415" />
                    <RANKING order="15" place="-1" resultid="13431" />
                    <RANKING order="16" place="-1" resultid="14310" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1118" agemax="12" agemin="12" name="12 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13197" />
                    <RANKING order="2" place="2" resultid="14550" />
                    <RANKING order="3" place="3" resultid="12452" />
                    <RANKING order="4" place="4" resultid="13711" />
                    <RANKING order="5" place="5" resultid="13215" />
                    <RANKING order="6" place="6" resultid="14613" />
                    <RANKING order="7" place="7" resultid="13227" />
                    <RANKING order="8" place="8" resultid="12353" />
                    <RANKING order="9" place="9" resultid="13655" />
                    <RANKING order="10" place="10" resultid="14120" />
                    <RANKING order="11" place="11" resultid="14531" />
                    <RANKING order="12" place="12" resultid="13534" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12936" daytime="11:22" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12937" daytime="11:24" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12938" daytime="11:26" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="12939" daytime="11:29" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="12940" daytime="11:31" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="12941" daytime="11:33" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="12942" daytime="11:35" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1119" daytime="11:37" gender="F" number="17" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <FEE currency="CHF" value="2000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1120" agemax="12" agemin="-1" name="12 Jahre und jünger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14651" />
                    <RANKING order="2" place="2" resultid="13553" />
                    <RANKING order="3" place="3" resultid="13555" />
                    <RANKING order="4" place="4" resultid="14652" />
                    <RANKING order="5" place="5" resultid="13740" />
                    <RANKING order="6" place="6" resultid="14666" />
                    <RANKING order="7" place="7" resultid="13204" />
                    <RANKING order="8" place="8" resultid="14347" />
                    <RANKING order="9" place="9" resultid="12461" />
                    <RANKING order="10" place="10" resultid="13742" />
                    <RANKING order="11" place="11" resultid="13206" />
                    <RANKING order="12" place="12" resultid="14349" />
                    <RANKING order="13" place="13" resultid="14350" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12944" daytime="11:37" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12945" daytime="11:41" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12946" daytime="11:45" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="14669" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1122" daytime="11:48" gender="M" number="18" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <FEE currency="CHF" value="2000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1123" agemax="12" agemin="-1" name="12 Jahre und jünger">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14650" />
                    <RANKING order="2" place="2" resultid="12457" />
                    <RANKING order="3" place="3" resultid="13202" />
                    <RANKING order="4" place="4" resultid="12459" />
                    <RANKING order="5" place="5" resultid="14345" />
                    <RANKING order="6" place="6" resultid="13738" />
                    <RANKING order="7" place="7" resultid="14665" />
                    <RANKING order="8" place="-1" resultid="13248" />
                    <RANKING order="9" place="-1" resultid="14346" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12947" daytime="11:48" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12948" daytime="11:52" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="14668" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
          <JUDGES>
            <JUDGE officialid="14677" role="REF" />
          </JUDGES>
        </SESSION>
        <SESSION date="2021-09-18" daytime="14:00" endtime="18:30" name="Nachmittag" number="2" officialmeeting="13:30" teamleadermeeting="13:15" warmupfrom="13:00" warmupuntil="13:45">
          <EVENTS>
            <EVENT eventid="1125" daytime="14:00" gender="F" number="19" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1128" agemax="14" agemin="13" name="13 und 14 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13474" />
                    <RANKING order="2" place="2" resultid="13669" />
                    <RANKING order="3" place="3" resultid="14587" />
                    <RANKING order="4" place="4" resultid="13641" />
                    <RANKING order="5" place="5" resultid="12368" />
                    <RANKING order="6" place="6" resultid="14607" />
                    <RANKING order="7" place="7" resultid="13184" />
                    <RANKING order="8" place="8" resultid="13087" />
                    <RANKING order="9" place="9" resultid="13705" />
                    <RANKING order="10" place="10" resultid="13720" />
                    <RANKING order="11" place="11" resultid="13485" />
                    <RANKING order="12" place="12" resultid="14603" />
                    <RANKING order="13" place="13" resultid="14540" />
                    <RANKING order="14" place="14" resultid="14231" />
                    <RANKING order="15" place="15" resultid="13117" />
                    <RANKING order="16" place="16" resultid="14619" />
                    <RANKING order="17" place="17" resultid="14595" />
                    <RANKING order="18" place="18" resultid="13052" />
                    <RANKING order="19" place="19" resultid="13136" />
                    <RANKING order="20" place="-1" resultid="13148" />
                    <RANKING order="21" place="-1" resultid="14050" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1129" agemax="16" agemin="15" name="15 und 16 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13047" />
                    <RANKING order="2" place="2" resultid="12377" />
                    <RANKING order="3" place="3" resultid="13687" />
                    <RANKING order="4" place="4" resultid="13716" />
                    <RANKING order="5" place="5" resultid="14647" />
                    <RANKING order="6" place="6" resultid="13142" />
                    <RANKING order="7" place="-1" resultid="13616" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1127" agemax="-1" agemin="17" name="17 und älter">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13702" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12949" daytime="14:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12950" daytime="14:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12951" daytime="14:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="12952" daytime="14:06" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="12953" daytime="14:08" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="12954" daytime="14:10" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="12955" daytime="14:12" number="7" order="7" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="*" timestandardlistid="5607">
                  <FEE currency="CHF" value="1000" />
                </TIMESTANDARDREF>
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1131" daytime="14:14" gender="M" number="20" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1132" agemax="14" agemin="13" name="13 und 14 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13637" />
                    <RANKING order="2" place="2" resultid="13158" />
                    <RANKING order="3" place="3" resultid="13168" />
                    <RANKING order="4" place="4" resultid="14333" />
                    <RANKING order="5" place="5" resultid="14579" />
                    <RANKING order="6" place="6" resultid="13111" />
                    <RANKING order="7" place="7" resultid="14174" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1133" agemax="16" agemin="15" name="15 und 16 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13519" />
                    <RANKING order="2" place="2" resultid="13072" />
                    <RANKING order="3" place="3" resultid="14631" />
                    <RANKING order="4" place="4" resultid="13608" />
                    <RANKING order="5" place="5" resultid="13795" />
                    <RANKING order="6" place="6" resultid="13174" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1135" agemax="-1" agemin="17" name="17 und älter">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13164" />
                    <RANKING order="2" place="2" resultid="12410" />
                    <RANKING order="3" place="3" resultid="13229" />
                    <RANKING order="4" place="-1" resultid="13066" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12957" daytime="14:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12958" daytime="14:16" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12959" daytime="14:18" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="12960" daytime="14:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="14653" daytime="14:21" number="5" order="5" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF marker="*" timestandardlistid="5605">
                  <FEE currency="CHF" value="1000" />
                </TIMESTANDARDREF>
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1136" daytime="14:24" gender="F" number="21" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1137" agemax="14" agemin="13" name="13 und 14 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14217" />
                    <RANKING order="2" place="2" resultid="14299" />
                    <RANKING order="3" place="3" resultid="13088" />
                    <RANKING order="4" place="4" resultid="13788" />
                    <RANKING order="5" place="5" resultid="13185" />
                    <RANKING order="6" place="6" resultid="14525" />
                    <RANKING order="7" place="7" resultid="14544" />
                    <RANKING order="8" place="8" resultid="12429" />
                    <RANKING order="9" place="9" resultid="13118" />
                    <RANKING order="10" place="10" resultid="13137" />
                    <RANKING order="11" place="11" resultid="14560" />
                    <RANKING order="12" place="12" resultid="13433" />
                    <RANKING order="13" place="13" resultid="14134" />
                    <RANKING order="14" place="14" resultid="13418" />
                    <RANKING order="15" place="15" resultid="13053" />
                    <RANKING order="16" place="16" resultid="12425" />
                    <RANKING order="17" place="17" resultid="14196" />
                    <RANKING order="18" place="-1" resultid="14158" />
                    <RANKING order="19" place="-1" resultid="13149" />
                    <RANKING order="20" place="-1" resultid="14055" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1138" agemax="16" agemin="15" name="15 und 16 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14672" />
                    <RANKING order="2" place="2" resultid="13516" />
                    <RANKING order="3" place="3" resultid="12376" />
                    <RANKING order="4" place="4" resultid="13540" />
                    <RANKING order="5" place="5" resultid="13717" />
                    <RANKING order="6" place="6" resultid="14249" />
                    <RANKING order="7" place="7" resultid="13143" />
                    <RANKING order="8" place="8" resultid="13440" />
                    <RANKING order="9" place="-1" resultid="13620" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1140" agemax="-1" agemin="17" name="17 und älter">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13612" />
                    <RANKING order="2" place="-1" resultid="13422" />
                    <RANKING order="3" place="-1" resultid="13509" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12962" daytime="14:24" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12963" daytime="14:26" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12964" daytime="14:29" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="12965" daytime="14:31" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="12966" daytime="14:33" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="12967" daytime="14:35" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="12968" daytime="14:37" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="12969" daytime="14:39" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1141" daytime="14:42" gender="M" number="22" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1142" agemax="14" agemin="13" name="13 und 14 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13792" />
                    <RANKING order="2" place="2" resultid="13728" />
                    <RANKING order="3" place="3" resultid="14567" />
                    <RANKING order="4" place="4" resultid="13169" />
                    <RANKING order="5" place="5" resultid="13523" />
                    <RANKING order="6" place="6" resultid="14334" />
                    <RANKING order="7" place="7" resultid="13159" />
                    <RANKING order="8" place="8" resultid="13543" />
                    <RANKING order="9" place="9" resultid="14629" />
                    <RANKING order="10" place="10" resultid="13625" />
                    <RANKING order="11" place="11" resultid="14552" />
                    <RANKING order="12" place="12" resultid="13112" />
                    <RANKING order="13" place="13" resultid="14599" />
                    <RANKING order="14" place="14" resultid="12433" />
                    <RANKING order="15" place="15" resultid="14191" />
                    <RANKING order="16" place="16" resultid="13428" />
                    <RANKING order="17" place="-1" resultid="13683" />
                    <RANKING order="18" place="-1" resultid="14623" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1143" agemax="16" agemin="15" name="15 und 16 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13499" />
                    <RANKING order="2" place="2" resultid="13073" />
                    <RANKING order="3" place="3" resultid="13785" />
                    <RANKING order="4" place="4" resultid="13782" />
                    <RANKING order="5" place="5" resultid="13175" />
                    <RANKING order="6" place="6" resultid="13778" />
                    <RANKING order="7" place="-1" resultid="14179" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1145" agemax="-1" agemin="17" name="17 und älter">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13245" />
                    <RANKING order="2" place="2" resultid="12372" />
                    <RANKING order="3" place="3" resultid="14258" />
                    <RANKING order="4" place="4" resultid="12338" />
                    <RANKING order="5" place="-1" resultid="13067" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12970" daytime="14:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12971" daytime="14:44" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12972" daytime="14:47" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="12973" daytime="14:49" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="12974" daytime="14:51" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="12975" daytime="14:53" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="12976" daytime="14:55" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="12977" daytime="14:57" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1146" daytime="14:59" gender="F" number="23" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1147" agemax="14" agemin="13" name="13 und 14 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13475" />
                    <RANKING order="2" place="2" resultid="13496" />
                    <RANKING order="3" place="3" resultid="12369" />
                    <RANKING order="4" place="4" resultid="13670" />
                    <RANKING order="5" place="5" resultid="14218" />
                    <RANKING order="6" place="6" resultid="14300" />
                    <RANKING order="7" place="7" resultid="13486" />
                    <RANKING order="8" place="8" resultid="13089" />
                    <RANKING order="9" place="9" resultid="13721" />
                    <RANKING order="10" place="10" resultid="14604" />
                    <RANKING order="11" place="11" resultid="14232" />
                    <RANKING order="12" place="12" resultid="14608" />
                    <RANKING order="13" place="13" resultid="14588" />
                    <RANKING order="14" place="14" resultid="14545" />
                    <RANKING order="15" place="15" resultid="14312" />
                    <RANKING order="16" place="16" resultid="13657" />
                    <RANKING order="17" place="17" resultid="14596" />
                    <RANKING order="18" place="18" resultid="14161" />
                    <RANKING order="19" place="19" resultid="13186" />
                    <RANKING order="20" place="20" resultid="14526" />
                    <RANKING order="21" place="21" resultid="13549" />
                    <RANKING order="22" place="22" resultid="14620" />
                    <RANKING order="23" place="23" resultid="13512" />
                    <RANKING order="24" place="24" resultid="13138" />
                    <RANKING order="25" place="25" resultid="13119" />
                    <RANKING order="26" place="26" resultid="13434" />
                    <RANKING order="27" place="27" resultid="14561" />
                    <RANKING order="28" place="28" resultid="13054" />
                    <RANKING order="29" place="29" resultid="13419" />
                    <RANKING order="30" place="30" resultid="14154" />
                    <RANKING order="31" place="31" resultid="14135" />
                    <RANKING order="32" place="32" resultid="12426" />
                    <RANKING order="33" place="-1" resultid="14541" />
                    <RANKING order="34" place="-1" resultid="13150" />
                    <RANKING order="35" place="-1" resultid="14052" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1148" agemax="16" agemin="15" name="15 und 16 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13463" />
                    <RANKING order="2" place="2" resultid="13048" />
                    <RANKING order="3" place="3" resultid="13507" />
                    <RANKING order="4" place="4" resultid="13645" />
                    <RANKING order="5" place="5" resultid="13199" />
                    <RANKING order="6" place="6" resultid="13688" />
                    <RANKING order="7" place="7" resultid="13629" />
                    <RANKING order="8" place="8" resultid="14250" />
                    <RANKING order="9" place="8" resultid="14643" />
                    <RANKING order="10" place="10" resultid="13517" />
                    <RANKING order="11" place="11" resultid="14648" />
                    <RANKING order="12" place="12" resultid="13144" />
                    <RANKING order="13" place="-1" resultid="13621" />
                    <RANKING order="14" place="-1" resultid="13617" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1150" agemax="-1" agemin="17" name="17 und älter">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13489" />
                    <RANKING order="2" place="2" resultid="14316" />
                    <RANKING order="3" place="3" resultid="13613" />
                    <RANKING order="4" place="4" resultid="13210" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12978" daytime="14:59" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12979" daytime="15:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12980" daytime="15:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="12981" daytime="15:06" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="12982" daytime="15:08" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="12983" daytime="15:10" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="12984" daytime="15:12" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="12985" daytime="15:14" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="12986" daytime="15:16" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="12987" daytime="15:17" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="12988" daytime="15:19" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="12989" daytime="15:21" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="12990" daytime="15:23" number="13" order="13" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1151" daytime="15:25" gender="M" number="24" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1152" agemax="14" agemin="13" name="13 und 14 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13713" />
                    <RANKING order="2" place="2" resultid="13729" />
                    <RANKING order="3" place="3" resultid="13638" />
                    <RANKING order="4" place="4" resultid="14568" />
                    <RANKING order="5" place="5" resultid="13170" />
                    <RANKING order="6" place="6" resultid="14335" />
                    <RANKING order="7" place="7" resultid="14580" />
                    <RANKING order="8" place="8" resultid="13160" />
                    <RANKING order="9" place="9" resultid="13530" />
                    <RANKING order="10" place="10" resultid="14175" />
                    <RANKING order="11" place="11" resultid="13113" />
                    <RANKING order="12" place="12" resultid="12421" />
                    <RANKING order="13" place="13" resultid="14600" />
                    <RANKING order="14" place="14" resultid="14192" />
                    <RANKING order="15" place="-1" resultid="14553" />
                    <RANKING order="16" place="-1" resultid="14624" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1153" agemax="16" agemin="15" name="15 und 16 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13074" />
                    <RANKING order="2" place="2" resultid="14288" />
                    <RANKING order="3" place="3" resultid="13695" />
                    <RANKING order="4" place="4" resultid="13520" />
                    <RANKING order="5" place="5" resultid="13176" />
                    <RANKING order="6" place="6" resultid="13796" />
                    <RANKING order="7" place="7" resultid="13609" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1155" agemax="-1" agemin="17" name="17 und älter">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12411" />
                    <RANKING order="2" place="2" resultid="14259" />
                    <RANKING order="3" place="3" resultid="13246" />
                    <RANKING order="4" place="4" resultid="13230" />
                    <RANKING order="5" place="5" resultid="14168" />
                    <RANKING order="6" place="-1" resultid="13068" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12991" daytime="15:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12992" daytime="15:27" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12993" daytime="15:29" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="12994" daytime="15:31" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="12995" daytime="15:33" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="12996" daytime="15:35" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="12997" daytime="15:37" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1156" daytime="15:39" gender="F" number="25" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1157" agemax="14" agemin="13" name="13 und 14 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14219" />
                    <RANKING order="2" place="2" resultid="14313" />
                    <RANKING order="3" place="3" resultid="13706" />
                    <RANKING order="4" place="4" resultid="13642" />
                    <RANKING order="5" place="5" resultid="14233" />
                    <RANKING order="6" place="6" resultid="14162" />
                    <RANKING order="7" place="7" resultid="12430" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1158" agemax="16" agemin="15" name="15 und 16 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13049" />
                    <RANKING order="2" place="2" resultid="13506" />
                    <RANKING order="3" place="3" resultid="13200" />
                    <RANKING order="4" place="4" resultid="14251" />
                    <RANKING order="5" place="5" resultid="14644" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1160" agemax="-1" agemin="17" name="17 und älter">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13703" />
                    <RANKING order="2" place="2" resultid="14317" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12998" daytime="15:39" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12999" daytime="15:43" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="13000" daytime="15:46" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="13001" daytime="15:49" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1161" daytime="15:52" gender="M" number="26" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1162" agemax="14" agemin="13" name="13 und 14 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13524" />
                    <RANKING order="2" place="2" resultid="14627" />
                    <RANKING order="3" place="3" resultid="13544" />
                    <RANKING order="4" place="4" resultid="14176" />
                    <RANKING order="5" place="5" resultid="12434" />
                    <RANKING order="6" place="6" resultid="14193" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1163" agemax="16" agemin="15" name="15 und 16 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14632" />
                    <RANKING order="2" place="2" resultid="13500" />
                    <RANKING order="3" place="3" resultid="14289" />
                    <RANKING order="4" place="-1" resultid="14180" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1165" agemax="-1" agemin="17" name="17 und älter">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13165" />
                    <RANKING order="2" place="2" resultid="12373" />
                    <RANKING order="3" place="3" resultid="12339" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="13003" daytime="15:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="13004" daytime="15:55" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="13005" daytime="15:59" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="13006" daytime="16:02" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1166" daytime="16:05" gender="F" number="27" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1167" agemax="14" agemin="13" name="13 und 14 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13671" />
                    <RANKING order="2" place="2" resultid="14301" />
                    <RANKING order="3" place="3" resultid="12370" />
                    <RANKING order="4" place="4" resultid="13487" />
                    <RANKING order="5" place="5" resultid="13789" />
                    <RANKING order="6" place="6" resultid="13658" />
                    <RANKING order="7" place="7" resultid="13090" />
                    <RANKING order="8" place="8" resultid="14159" />
                    <RANKING order="9" place="9" resultid="13120" />
                    <RANKING order="10" place="10" resultid="13055" />
                    <RANKING order="11" place="11" resultid="13139" />
                    <RANKING order="12" place="12" resultid="12427" />
                    <RANKING order="13" place="13" resultid="13513" />
                    <RANKING order="14" place="14" resultid="13550" />
                    <RANKING order="15" place="15" resultid="14156" />
                    <RANKING order="16" place="16" resultid="14136" />
                    <RANKING order="17" place="17" resultid="14197" />
                    <RANKING order="18" place="-1" resultid="13151" />
                    <RANKING order="19" place="-1" resultid="14051" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1168" agemax="16" agemin="15" name="15 und 16 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14671" />
                    <RANKING order="2" place="2" resultid="13464" />
                    <RANKING order="3" place="3" resultid="13646" />
                    <RANKING order="4" place="4" resultid="13145" />
                    <RANKING order="5" place="-1" resultid="13622" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1170" agemax="-1" agemin="17" name="17 und älter">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13490" />
                    <RANKING order="2" place="2" resultid="13614" />
                    <RANKING order="3" place="-1" resultid="13510" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="13007" daytime="16:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="13008" daytime="16:07" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="13009" daytime="16:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="13010" daytime="16:12" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="13011" daytime="16:14" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="13012" daytime="16:16" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="14115" daytime="16:18" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1171" daytime="16:20" gender="M" number="28" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1172" agemax="14" agemin="13" name="13 und 14 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13714" />
                    <RANKING order="2" place="2" resultid="13639" />
                    <RANKING order="3" place="3" resultid="13171" />
                    <RANKING order="4" place="4" resultid="14336" />
                    <RANKING order="5" place="5" resultid="13161" />
                    <RANKING order="6" place="6" resultid="12422" />
                    <RANKING order="7" place="7" resultid="13114" />
                    <RANKING order="8" place="8" resultid="13626" />
                    <RANKING order="9" place="9" resultid="13684" />
                    <RANKING order="10" place="-1" resultid="13793" />
                    <RANKING order="11" place="-1" resultid="14625" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1173" agemax="16" agemin="15" name="15 und 16 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13075" />
                    <RANKING order="2" place="2" resultid="13696" />
                    <RANKING order="3" place="3" resultid="13786" />
                    <RANKING order="4" place="4" resultid="13783" />
                    <RANKING order="5" place="5" resultid="13177" />
                    <RANKING order="6" place="6" resultid="13779" />
                    <RANKING order="7" place="-1" resultid="14181" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1175" agemax="-1" agemin="17" name="17 und älter">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12409" />
                    <RANKING order="2" place="2" resultid="14260" />
                    <RANKING order="3" place="3" resultid="14169" />
                    <RANKING order="4" place="-1" resultid="13069" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="13013" daytime="16:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="13014" daytime="16:23" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="13015" daytime="16:25" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="13016" daytime="16:27" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="13017" daytime="16:29" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="13018" daytime="16:31" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1176" daytime="16:33" gender="F" number="29" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1177" agemax="14" agemin="13" name="13 und 14 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13497" />
                    <RANKING order="2" place="2" resultid="14220" />
                    <RANKING order="3" place="3" resultid="13722" />
                    <RANKING order="4" place="4" resultid="13091" />
                    <RANKING order="5" place="5" resultid="14302" />
                    <RANKING order="6" place="6" resultid="14546" />
                    <RANKING order="7" place="7" resultid="14605" />
                    <RANKING order="8" place="8" resultid="14314" />
                    <RANKING order="9" place="9" resultid="14609" />
                    <RANKING order="10" place="10" resultid="14597" />
                    <RANKING order="11" place="11" resultid="13643" />
                    <RANKING order="12" place="12" resultid="13707" />
                    <RANKING order="13" place="13" resultid="14589" />
                    <RANKING order="14" place="14" resultid="14160" />
                    <RANKING order="15" place="15" resultid="14234" />
                    <RANKING order="16" place="16" resultid="13790" />
                    <RANKING order="17" place="17" resultid="13659" />
                    <RANKING order="18" place="18" resultid="13187" />
                    <RANKING order="19" place="19" resultid="14527" />
                    <RANKING order="20" place="20" resultid="14542" />
                    <RANKING order="21" place="21" resultid="13551" />
                    <RANKING order="22" place="22" resultid="14621" />
                    <RANKING order="23" place="23" resultid="13140" />
                    <RANKING order="24" place="24" resultid="12431" />
                    <RANKING order="25" place="25" resultid="13121" />
                    <RANKING order="26" place="26" resultid="13514" />
                    <RANKING order="27" place="27" resultid="13435" />
                    <RANKING order="28" place="28" resultid="13420" />
                    <RANKING order="29" place="29" resultid="14562" />
                    <RANKING order="30" place="30" resultid="14137" />
                    <RANKING order="31" place="31" resultid="13056" />
                    <RANKING order="32" place="32" resultid="14155" />
                    <RANKING order="33" place="33" resultid="14198" />
                    <RANKING order="34" place="-1" resultid="13152" />
                    <RANKING order="35" place="-1" resultid="14054" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1178" agemax="16" agemin="15" name="15 und 16 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13050" />
                    <RANKING order="2" place="2" resultid="13541" />
                    <RANKING order="3" place="3" resultid="12378" />
                    <RANKING order="4" place="4" resultid="13201" />
                    <RANKING order="5" place="5" resultid="13689" />
                    <RANKING order="6" place="6" resultid="13647" />
                    <RANKING order="7" place="7" resultid="14645" />
                    <RANKING order="8" place="8" resultid="14252" />
                    <RANKING order="9" place="9" resultid="13718" />
                    <RANKING order="10" place="10" resultid="13146" />
                    <RANKING order="11" place="11" resultid="14649" />
                    <RANKING order="12" place="12" resultid="13441" />
                    <RANKING order="13" place="-1" resultid="13623" />
                    <RANKING order="14" place="-1" resultid="13618" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1180" agemax="-1" agemin="17" name="17 und älter">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14318" />
                    <RANKING order="2" place="2" resultid="13211" />
                    <RANKING order="3" place="3" resultid="13423" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="13019" daytime="16:33" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="13020" daytime="16:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="13021" daytime="16:37" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="13022" daytime="16:39" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="13023" daytime="16:41" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="13024" daytime="16:43" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="13025" daytime="16:44" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="13026" daytime="16:46" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="13027" daytime="16:48" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="13028" daytime="16:49" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="13029" daytime="16:51" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="13030" daytime="16:53" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="13031" daytime="16:54" number="13" order="13" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1181" daytime="16:56" gender="M" number="30" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="CHF" value="1000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1182" agemax="14" agemin="13" name="13 und 14 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13730" />
                    <RANKING order="2" place="2" resultid="14569" />
                    <RANKING order="3" place="3" resultid="13172" />
                    <RANKING order="4" place="4" resultid="13162" />
                    <RANKING order="5" place="5" resultid="13115" />
                    <RANKING order="6" place="6" resultid="14177" />
                    <RANKING order="7" place="7" resultid="14628" />
                    <RANKING order="8" place="8" resultid="14581" />
                    <RANKING order="9" place="9" resultid="13685" />
                    <RANKING order="10" place="10" resultid="14554" />
                    <RANKING order="11" place="11" resultid="12423" />
                    <RANKING order="12" place="12" resultid="13627" />
                    <RANKING order="13" place="13" resultid="13531" />
                    <RANKING order="14" place="14" resultid="12435" />
                    <RANKING order="15" place="15" resultid="14601" />
                    <RANKING order="16" place="16" resultid="14194" />
                    <RANKING order="17" place="17" resultid="13429" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1183" agemax="16" agemin="15" name="15 und 16 Jahre">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="14290" />
                    <RANKING order="2" place="2" resultid="14633" />
                    <RANKING order="3" place="3" resultid="13610" />
                    <RANKING order="4" place="4" resultid="13076" />
                    <RANKING order="5" place="5" resultid="13521" />
                    <RANKING order="6" place="6" resultid="13178" />
                    <RANKING order="7" place="7" resultid="13780" />
                    <RANKING order="8" place="-1" resultid="14182" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1185" agemax="-1" agemin="17" name="17 und älter">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13166" />
                    <RANKING order="2" place="2" resultid="12374" />
                    <RANKING order="3" place="3" resultid="14261" />
                    <RANKING order="4" place="4" resultid="13247" />
                    <RANKING order="5" place="5" resultid="12340" />
                    <RANKING order="6" place="6" resultid="13231" />
                    <RANKING order="7" place="7" resultid="14170" />
                    <RANKING order="8" place="-1" resultid="13070" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="13033" daytime="16:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="13034" daytime="16:58" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="13035" daytime="17:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="13036" daytime="17:02" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="13037" daytime="17:04" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="13038" daytime="17:05" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="13039" daytime="17:07" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="13040" daytime="17:08" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="14655" daytime="17:10" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1186" daytime="17:12" gender="F" number="31" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="CHF" value="2000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1190" agemax="-1" agemin="13" name="13 und älter">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13554" />
                    <RANKING order="2" place="2" resultid="13741" />
                    <RANKING order="3" place="3" resultid="13556" />
                    <RANKING order="4" place="4" resultid="13743" />
                    <RANKING order="5" place="5" resultid="13205" />
                    <RANKING order="6" place="6" resultid="14348" />
                    <RANKING order="7" place="7" resultid="12460" />
                    <RANKING order="8" place="8" resultid="13207" />
                    <RANKING order="9" place="9" resultid="13445" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="13041" daytime="17:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="13042" daytime="17:18" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="13043" daytime="17:23" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1191" daytime="17:28" gender="M" number="32" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="CHF" value="2000" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1192" agemax="-1" agemin="13" name="13 und älter">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="13739" />
                    <RANKING order="2" place="2" resultid="13203" />
                    <RANKING order="3" place="3" resultid="13797" />
                    <RANKING order="4" place="4" resultid="12458" />
                    <RANKING order="5" place="5" resultid="13552" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="13044" daytime="17:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="13045" daytime="17:33" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
          <JUDGES>
            <JUDGE officialid="14677" role="REF" />
          </JUDGES>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="FTAL" nation="SUI" region="RZW" clubid="12480" name="Schwimmclub Fricktal">
          <ATHLETES>
            <ATHLETE firstname="Jael" lastname="Schweizer" birthdate="2012-11-08" gender="F" nation="SUI" athleteid="14291">
              <RESULTS>
                <RESULT eventid="1073" points="77" swimtime="00:01:00.08" resultid="14292" heatid="12872" lane="2" entrytime="00:00:59.45" entrycourse="LCM" />
                <RESULT eventid="1092" points="103" swimtime="00:01:00.82" resultid="14293" heatid="12887" lane="1" entrytime="00:01:09.01" entrycourse="LCM" />
                <RESULT eventid="1106" points="81" swimtime="00:00:52.93" resultid="14294" heatid="12913" lane="3" entrytime="00:00:55.94" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joshua" lastname="Weibel" birthdate="2007-03-15" gender="M" nation="SUI" license="112081" athleteid="14332">
              <RESULTS>
                <RESULT eventid="1131" points="217" swimtime="00:01:19.51" resultid="14333" heatid="12958" lane="2" entrytime="00:01:20.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="250" swimtime="00:01:16.66" resultid="14334" heatid="12974" lane="1" entrytime="00:01:20.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="257" swimtime="00:01:17.49" resultid="14335" heatid="12992" lane="4" entrytime="00:01:34.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="239" swimtime="00:01:29.14" resultid="14336" heatid="13014" lane="1" entrytime="00:01:44.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carina" lastname="Sutter" birthdate="2007-04-16" gender="F" nation="SUI" license="109162" athleteid="14311">
              <RESULTS>
                <RESULT eventid="1146" points="349" swimtime="00:01:20.26" resultid="14312" heatid="12983" lane="1" entrytime="00:01:24.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="444" swimtime="00:02:24.73" resultid="14313" heatid="12999" lane="3" entrytime="00:02:32.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.88" />
                    <SPLIT distance="100" swimtime="00:01:09.84" />
                    <SPLIT distance="150" swimtime="00:01:48.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="398" swimtime="00:01:08.28" resultid="14314" heatid="13025" lane="4" entrytime="00:01:09.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Linda" lastname="Egger" birthdate="2007-08-15" gender="F" nation="SUI" license="109159" athleteid="14216">
              <RESULTS>
                <RESULT eventid="1136" points="467" swimtime="00:01:10.73" resultid="14217" heatid="12968" lane="4" entrytime="00:01:14.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="428" swimtime="00:01:14.98" resultid="14218" heatid="12987" lane="3" entrytime="00:01:18.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="453" swimtime="00:02:23.74" resultid="14219" heatid="13000" lane="1" entrytime="00:02:26.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.58" />
                    <SPLIT distance="100" swimtime="00:01:08.38" />
                    <SPLIT distance="150" swimtime="00:01:45.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="473" swimtime="00:01:04.48" resultid="14220" heatid="13029" lane="1" entrytime="00:01:05.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nela" lastname="Hanak" birthdate="2012-04-12" gender="F" nation="SUI" license="122842" athleteid="14253">
              <RESULTS>
                <RESULT eventid="1073" points="130" swimtime="00:00:50.51" resultid="14254" heatid="12876" lane="4" entrytime="00:00:53.91" entrycourse="LCM" />
                <RESULT eventid="1092" points="162" swimtime="00:00:52.33" resultid="14255" heatid="14113" lane="3" entrytime="00:00:52.72" entrycourse="LCM" />
                <RESULT eventid="1106" points="98" swimtime="00:00:49.72" resultid="14256" heatid="12917" lane="4" entrytime="00:00:46.73" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Noa" lastname="Sutter" birthdate="2010-08-05" gender="M" nation="SUI" license="119865" athleteid="14319">
              <RESULTS>
                <RESULT comment="504 - Brustbeinschlag während des Schwimmens" eventid="1060" status="DSQ" swimtime="00:00:55.25" resultid="14320" heatid="12852" lane="3" entrytime="00:00:56.00" />
                <RESULT eventid="1103" points="123" swimtime="00:01:51.18" resultid="14321" heatid="12907" lane="2" entrytime="00:02:00.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="59" swimtime="00:01:55.19" resultid="14322" heatid="12938" lane="4" entrytime="00:01:43.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1070" points="72" swimtime="00:01:56.11" resultid="14323" heatid="12865" lane="1" entrytime="00:01:57.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leon" lastname="Shala" birthdate="2011-03-03" gender="M" nation="SUI" athleteid="14295">
              <RESULTS>
                <RESULT comment="306 - Wand in Bauchlage verlassen  (Wende ...)" eventid="1076" status="DSQ" swimtime="00:01:06.25" resultid="14296" heatid="12880" lane="2" entrytime="00:01:00.00" />
                <RESULT eventid="1109" points="38" swimtime="00:00:59.57" resultid="14297" heatid="12920" lane="3" entrytime="00:00:56.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arik" lastname="Benz" birthdate="2012-06-05" gender="M" nation="SUI" athleteid="14207">
              <RESULTS>
                <RESULT eventid="1060" points="62" swimtime="00:00:54.83" resultid="14208" heatid="12854" lane="4" entrytime="00:00:49.44" entrycourse="LCM" />
                <RESULT eventid="1076" points="80" swimtime="00:00:51.51" resultid="14209" heatid="12881" lane="1" entrytime="00:00:57.26" entrycourse="LCM" />
                <RESULT eventid="1096" points="60" swimtime="00:01:04.35" resultid="14210" heatid="12893" lane="2" entrytime="00:01:02.66" entrycourse="LCM" />
                <RESULT eventid="1109" points="121" swimtime="00:00:40.71" resultid="14211" heatid="12923" lane="1" entrytime="00:00:41.29" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amélie" lastname="Friesewinkel" birthdate="2011-02-04" gender="F" nation="SUI" athleteid="14225">
              <RESULTS>
                <RESULT eventid="1073" points="109" swimtime="00:00:53.51" resultid="14226" heatid="12876" lane="1" entrytime="00:00:53.59" entrycourse="LCM" />
                <RESULT eventid="1092" points="129" swimtime="00:00:56.47" resultid="14227" heatid="12890" lane="1" entrytime="00:00:59.05" entrycourse="LCM" />
                <RESULT eventid="1106" points="131" swimtime="00:00:45.09" resultid="14228" heatid="12917" lane="1" entrytime="00:00:45.88" entrycourse="LCM" />
                <RESULT eventid="1053" points="66" swimtime="00:01:00.25" resultid="14229" heatid="12846" lane="2" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lena" lastname="Nikolic" birthdate="2012-01-01" gender="F" nation="SUI" athleteid="14283">
              <RESULTS>
                <RESULT comment="302 - Wand nicht berührt (Wende ...)" eventid="1073" status="DSQ" swimtime="00:00:52.28" resultid="14284" heatid="12874" lane="3" entrytime="00:00:55.00" />
                <RESULT eventid="1092" points="56" swimtime="00:01:14.47" resultid="14285" heatid="12888" lane="4" entrytime="00:01:05.00" />
                <RESULT eventid="1106" points="77" swimtime="00:00:53.87" resultid="14286" heatid="12914" lane="1" entrytime="00:00:51.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Soraya" lastname="Euler" birthdate="2013-03-29" gender="F" nation="SUI" athleteid="14221">
              <RESULTS>
                <RESULT eventid="1073" points="28" swimtime="00:01:23.64" resultid="14222" heatid="12870" lane="3" />
                <RESULT eventid="1092" points="52" swimtime="00:01:16.10" resultid="14223" heatid="12886" lane="1" />
                <RESULT eventid="1106" points="16" swimtime="00:01:30.41" resultid="14224" heatid="12911" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juliette" lastname="Siegfried" birthdate="2008-04-11" gender="F" nation="SUI" license="109161" athleteid="14298">
              <RESULTS>
                <RESULT eventid="1136" points="415" swimtime="00:01:13.53" resultid="14299" heatid="12967" lane="3" entrytime="00:01:18.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="417" swimtime="00:01:15.60" resultid="14300" heatid="12986" lane="3" entrytime="00:01:19.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1166" points="420" swimtime="00:01:23.22" resultid="14301" heatid="13012" lane="3" entrytime="00:01:23.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="405" swimtime="00:01:07.87" resultid="14302" heatid="13025" lane="3" entrytime="00:01:09.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Selina" lastname="Unternaehrer" birthdate="2012-11-21" gender="F" nation="SUI" athleteid="14328">
              <RESULTS>
                <RESULT eventid="1073" points="68" swimtime="00:01:02.65" resultid="14329" heatid="12870" lane="1" />
                <RESULT eventid="1092" points="83" swimtime="00:01:05.40" resultid="14330" heatid="12885" lane="2" />
                <RESULT eventid="1106" points="55" swimtime="00:00:59.95" resultid="14331" heatid="12912" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Krzeminska" birthdate="2011-04-28" gender="F" nation="POL" athleteid="14271">
              <RESULTS>
                <RESULT comment="404 - Nicht in Rückenlage angeschlagen (Ziel)" eventid="1073" status="DSQ" swimtime="00:01:06.19" resultid="14272" heatid="12871" lane="1" />
                <RESULT comment="403 - Nicht mit beiden Händen gleichzeitig angeschlagen (Ziel)" eventid="1092" status="DSQ" swimtime="00:01:31.76" resultid="14273" heatid="12886" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nina" lastname="Wüthrich" birthdate="2012-11-25" gender="F" nation="SUI" license="122841" athleteid="14337">
              <RESULTS>
                <RESULT comment="304 - Schwimmen in Bauchlage vor der Wende (Wende ...)" eventid="1073" status="DSQ" swimtime="00:00:54.79" resultid="14338" heatid="12873" lane="2" entrytime="00:00:55.27" entrycourse="LCM" />
                <RESULT eventid="1092" points="139" swimtime="00:00:55.07" resultid="14339" heatid="12891" lane="3" entrytime="00:00:56.90" entrycourse="LCM" />
                <RESULT eventid="1106" points="77" swimtime="00:00:53.79" resultid="14340" heatid="12913" lane="2" entrytime="00:00:54.02" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elina" lastname="Gallert" birthdate="2007-05-12" gender="F" nation="SUI" license="107434" athleteid="14230">
              <RESULTS>
                <RESULT eventid="1125" points="292" swimtime="00:01:22.23" resultid="14231" heatid="12951" lane="1" entrytime="00:01:25.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="362" swimtime="00:01:19.24" resultid="14232" heatid="12984" lane="1" entrytime="00:01:23.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="387" swimtime="00:02:31.53" resultid="14233" heatid="12998" lane="2" entrytime="00:02:36.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.23" />
                    <SPLIT distance="100" swimtime="00:01:12.61" />
                    <SPLIT distance="150" swimtime="00:01:52.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="363" swimtime="00:01:10.41" resultid="14234" heatid="13023" lane="3" entrytime="00:01:11.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Xenia" lastname="Zolliker" birthdate="2010-10-19" gender="F" nation="SUI" license="119028" athleteid="14341">
              <RESULTS>
                <RESULT eventid="1053" points="97" swimtime="00:00:53.05" resultid="14342" heatid="12847" lane="1" entrytime="00:00:54.19" entrycourse="SCM" />
                <RESULT eventid="1084" points="173" swimtime="00:03:17.99" resultid="14343" heatid="12883" lane="3" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.10" />
                    <SPLIT distance="100" swimtime="00:01:34.82" />
                    <SPLIT distance="150" swimtime="00:02:28.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="155" swimtime="00:01:33.44" resultid="14344" heatid="12928" lane="2" entrytime="00:01:29.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Debora" lastname="Mettler" birthdate="2011-05-06" gender="F" nation="SUI" license="121723" athleteid="14278">
              <RESULTS>
                <RESULT eventid="1053" status="WDR" swimtime="00:00:00.00" resultid="14279" heatid="12846" lane="1" entrytime="00:00:55.00" />
                <RESULT eventid="1073" status="WDR" swimtime="00:00:00.00" resultid="14280" heatid="12874" lane="2" entrytime="00:00:54.87" entrycourse="LCM" />
                <RESULT eventid="1092" status="WDR" swimtime="00:00:00.00" resultid="14281" heatid="12889" lane="4" entrytime="00:01:00.01" entrycourse="LCM" />
                <RESULT eventid="1106" status="WDR" swimtime="00:00:00.00" resultid="14282" heatid="12915" lane="1" entrytime="00:00:48.68" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Loïc" lastname="Siegfried" birthdate="2012-10-16" gender="M" nation="SUI" license="122840" athleteid="14303">
              <RESULTS>
                <RESULT eventid="1060" points="71" swimtime="00:00:52.46" resultid="14304" heatid="12852" lane="2" entrytime="00:00:55.00" />
                <RESULT eventid="1076" points="86" swimtime="00:00:50.26" resultid="14305" heatid="12882" lane="2" entrytime="00:00:48.02" entrycourse="LCM" />
                <RESULT eventid="1096" points="89" swimtime="00:00:56.51" resultid="14306" heatid="12894" lane="3" entrytime="00:00:57.37" entrycourse="LCM" />
                <RESULT eventid="1109" points="93" swimtime="00:00:44.40" resultid="14307" heatid="12922" lane="2" entrytime="00:00:42.76" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mia" lastname="Gisler" birthdate="2006-07-29" gender="F" nation="SUI" license="116851" athleteid="14248">
              <RESULTS>
                <RESULT eventid="1136" points="354" swimtime="00:01:17.54" resultid="14249" heatid="12966" lane="4" entrytime="00:01:23.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="383" swimtime="00:01:17.80" resultid="14250" heatid="12983" lane="4" entrytime="00:01:24.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="437" swimtime="00:02:25.49" resultid="14251" heatid="12999" lane="2" entrytime="00:02:31.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.65" />
                    <SPLIT distance="100" swimtime="00:01:08.35" />
                    <SPLIT distance="150" swimtime="00:01:47.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="417" swimtime="00:01:07.26" resultid="14252" heatid="13024" lane="2" entrytime="00:01:09.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lewis" lastname="Rippstein" birthdate="2006-01-02" gender="M" nation="SUI" license="103726" athleteid="14287">
              <RESULTS>
                <RESULT eventid="1151" points="360" swimtime="00:01:09.24" resultid="14288" heatid="12995" lane="4" entrytime="00:01:18.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1161" points="354" swimtime="00:02:20.35" resultid="14289" heatid="13006" lane="4" entrytime="00:02:23.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.43" />
                    <SPLIT distance="100" swimtime="00:01:05.89" />
                    <SPLIT distance="150" swimtime="00:01:43.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="399" swimtime="00:01:01.04" resultid="14290" heatid="13040" lane="1" entrytime="00:01:01.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Larissa" lastname="Sutter" birthdate="2004-12-20" gender="F" nation="SUI" license="100332" athleteid="14315">
              <RESULTS>
                <RESULT eventid="1146" points="399" swimtime="00:01:16.72" resultid="14316" heatid="12988" lane="1" entrytime="00:01:17.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="434" swimtime="00:02:25.79" resultid="14317" heatid="13000" lane="2" entrytime="00:02:24.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.47" />
                    <SPLIT distance="100" swimtime="00:01:08.27" />
                    <SPLIT distance="150" swimtime="00:01:46.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="431" swimtime="00:01:06.49" resultid="14318" heatid="13030" lane="3" entrytime="00:01:04.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eric Keizo" lastname="Tomita" birthdate="2012-05-01" gender="M" nation="GER" athleteid="14324">
              <RESULTS>
                <RESULT eventid="1076" points="67" swimtime="00:00:54.58" resultid="14325" heatid="12880" lane="4" entrytime="00:01:03.99" entrycourse="LCM" />
                <RESULT eventid="1096" points="56" swimtime="00:01:05.91" resultid="14326" heatid="12893" lane="1" entrytime="00:01:05.38" entrycourse="LCM" />
                <RESULT eventid="1109" points="79" swimtime="00:00:46.94" resultid="14327" heatid="12921" lane="1" entrytime="00:00:49.84" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julius" lastname="Ilten" birthdate="2004-01-23" gender="M" nation="GER" license="106861" athleteid="14257">
              <RESULTS>
                <RESULT eventid="1141" points="360" swimtime="00:01:07.90" resultid="14258" heatid="12977" lane="3" entrytime="00:01:07.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="428" swimtime="00:01:05.39" resultid="14259" heatid="12997" lane="2" entrytime="00:01:06.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="410" swimtime="00:01:14.45" resultid="14260" heatid="13018" lane="4" entrytime="00:01:16.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="483" swimtime="00:00:57.24" resultid="14261" heatid="14655" lane="1" entrytime="00:00:57.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Liz" lastname="Geissler" birthdate="2010-10-23" gender="F" nation="SUI" athleteid="14239">
              <RESULTS>
                <RESULT eventid="1065" points="107" swimtime="00:01:55.34" resultid="14240" heatid="12857" lane="2" entrytime="00:01:54.24" entrycourse="LCM" />
                <RESULT eventid="1099" points="88" swimtime="00:02:19.80" resultid="14241" heatid="12897" lane="1" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="100" swimtime="00:01:47.96" resultid="14242" heatid="12926" lane="3" entrytime="00:01:46.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1053" points="46" swimtime="00:01:07.82" resultid="14243" heatid="12846" lane="3" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Raya" lastname="Benz" birthdate="2014-03-05" gender="F" nation="SUI" athleteid="14212">
              <RESULTS>
                <RESULT comment="404 - Nicht in Rückenlage angeschlagen (Ziel)" eventid="1073" status="DSQ" swimtime="00:01:21.33" resultid="14213" heatid="12870" lane="2" />
                <RESULT comment="521 - Körper nicht in Brustlage" eventid="1092" status="DSQ" swimtime="00:01:37.22" resultid="14214" heatid="12885" lane="1" />
                <RESULT eventid="1106" points="10" swimtime="00:01:44.41" resultid="14215" heatid="12911" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Noelle" lastname="Giess" birthdate="2012-02-16" gender="F" nation="SUI" athleteid="14244">
              <RESULTS>
                <RESULT comment="404 - Nicht in Rückenlage angeschlagen (Ziel)" eventid="1073" status="DSQ" swimtime="00:01:02.91" resultid="14245" heatid="12871" lane="4" />
                <RESULT comment="403 - Nicht mit beiden Händen gleichzeitig angeschlagen (Ziel)" eventid="1092" status="DSQ" swimtime="00:01:20.14" resultid="14246" heatid="12885" lane="3" />
                <RESULT eventid="1106" points="37" swimtime="00:01:08.71" resultid="14247" heatid="12911" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Norina" lastname="Gallert" birthdate="2011-12-11" gender="F" nation="SUI" license="121348" athleteid="14235">
              <RESULTS>
                <RESULT eventid="1073" points="129" swimtime="00:00:50.58" resultid="14236" heatid="12875" lane="2" entrytime="00:00:53.99" entrycourse="LCM" />
                <RESULT eventid="1092" points="133" swimtime="00:00:55.93" resultid="14237" heatid="12891" lane="2" entrytime="00:00:55.99" entrycourse="LCM" />
                <RESULT eventid="1106" points="111" swimtime="00:00:47.65" resultid="14238" heatid="12915" lane="4" entrytime="00:00:49.11" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theodor" lastname="Karotki" birthdate="2010-10-25" gender="M" nation="SUI" license="122766" athleteid="14262">
              <RESULTS>
                <RESULT eventid="1060" points="39" swimtime="00:01:04.12" resultid="14263" heatid="12852" lane="1" entrytime="00:00:58.00" />
                <RESULT eventid="1088" points="102" swimtime="00:03:32.51" resultid="14264" heatid="12884" lane="1" entrytime="00:03:08.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.38" />
                    <SPLIT distance="100" swimtime="00:01:40.52" />
                    <SPLIT distance="150" swimtime="00:02:37.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="107" swimtime="00:01:56.52" resultid="14265" heatid="12907" lane="4" entrytime="00:02:00.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="89" swimtime="00:01:40.64" resultid="14266" heatid="12938" lane="3" entrytime="00:01:35.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Konstantin" lastname="Stikhin" birthdate="2010-12-14" gender="M" nation="SUI" athleteid="14308">
              <RESULTS>
                <RESULT comment="304 - Schwimmen in Bauchlage vor der Wende (Wende ...)" eventid="1070" status="DSQ" swimtime="00:02:31.56" resultid="14309" heatid="12864" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" status="WDR" swimtime="00:00:00.00" resultid="14310" heatid="12936" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre" lastname="Kovac" birthdate="2012-08-02" gender="M" nation="SUI" athleteid="14267">
              <RESULTS>
                <RESULT comment="304 - Schwimmen in Bauchlage vor der Wende (Wende ...)" eventid="1076" status="DSQ" swimtime="00:01:15.34" resultid="14268" heatid="12878" lane="3" />
                <RESULT comment="526 - Beinbewegung nicht gleichzeitig in derselben horizontalen Ebene" eventid="1096" status="DSQ" swimtime="00:01:32.66" resultid="14269" heatid="12892" lane="1" />
                <RESULT eventid="1109" points="11" swimtime="00:01:29.99" resultid="14270" heatid="12919" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorine" lastname="Martin" birthdate="2009-04-26" gender="F" nation="SUI" athleteid="14274">
              <RESULTS>
                <RESULT eventid="1053" points="226" swimtime="00:00:40.01" resultid="14275" heatid="12851" lane="4" entrytime="00:00:40.00" />
                <RESULT eventid="1065" points="201" swimtime="00:01:33.63" resultid="14276" heatid="12861" lane="1" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="263" swimtime="00:01:18.41" resultid="14277" heatid="12932" lane="2" entrytime="00:01:21.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1122" points="94" swimtime="00:02:59.67" resultid="14345" heatid="12947" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.75" />
                    <SPLIT distance="100" swimtime="00:01:30.91" />
                    <SPLIT distance="150" swimtime="00:02:12.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14262" number="1" />
                    <RELAYPOSITION athleteid="14319" number="2" />
                    <RELAYPOSITION athleteid="14207" number="3" />
                    <RELAYPOSITION athleteid="14303" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1191" points="366" status="EXH" swimtime="00:04:15.85" resultid="14675" heatid="13044" lane="1">
                  <SPLITS>
                    <SPLIT distance="300" swimtime="00:03:15.53" />
                    <SPLIT distance="350" swimtime="00:03:44.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14257" number="1" />
                    <RELAYPOSITION athleteid="13157" number="2" />
                    <RELAYPOSITION athleteid="14332" number="3" />
                    <RELAYPOSITION athleteid="14287" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT comment="302 - Wand nicht berührt (Wende 3)" eventid="1122" status="DSQ" swimtime="00:03:59.66" resultid="14346" heatid="12947" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.30" />
                    <SPLIT distance="100" swimtime="00:01:47.49" />
                    <SPLIT distance="150" swimtime="00:03:14.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14324" number="1" />
                    <RELAYPOSITION athleteid="14295" number="2" />
                    <RELAYPOSITION athleteid="14267" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="13077" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1119" points="172" swimtime="00:02:46.30" resultid="14347" heatid="12944" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.86" />
                    <SPLIT distance="100" swimtime="00:01:18.82" />
                    <SPLIT distance="150" swimtime="00:02:03.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14274" number="1" />
                    <RELAYPOSITION athleteid="14341" number="2" />
                    <RELAYPOSITION athleteid="14253" number="3" />
                    <RELAYPOSITION athleteid="14225" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1186" points="433" swimtime="00:04:32.95" resultid="14348" heatid="13041" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.74" />
                    <SPLIT distance="100" swimtime="00:01:08.62" />
                    <SPLIT distance="150" swimtime="00:01:40.32" />
                    <SPLIT distance="200" swimtime="00:02:17.83" />
                    <SPLIT distance="250" swimtime="00:02:50.99" />
                    <SPLIT distance="300" swimtime="00:03:27.06" />
                    <SPLIT distance="350" swimtime="00:03:57.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14315" number="1" />
                    <RELAYPOSITION athleteid="14298" number="2" />
                    <RELAYPOSITION athleteid="14311" number="3" />
                    <RELAYPOSITION athleteid="14216" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1119" points="96" swimtime="00:03:21.41" resultid="14349" heatid="12944" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.26" />
                    <SPLIT distance="100" swimtime="00:01:40.69" />
                    <SPLIT distance="150" swimtime="00:02:33.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14239" number="1" />
                    <RELAYPOSITION athleteid="14337" number="2" />
                    <RELAYPOSITION athleteid="14283" number="3" />
                    <RELAYPOSITION athleteid="14235" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="3">
              <RESULTS>
                <RESULT eventid="1119" points="41" swimtime="00:04:28.01" resultid="14350" heatid="12945" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.99" />
                    <SPLIT distance="100" swimtime="00:01:53.29" />
                    <SPLIT distance="150" swimtime="00:02:59.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14291" number="1" />
                    <RELAYPOSITION athleteid="14328" number="2" />
                    <RELAYPOSITION athleteid="14244" number="3" />
                    <RELAYPOSITION athleteid="14221" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
          <COACHES>
            <COACH firstname="Agnieszka" gender="F" lastname="Bujoczek" nation="POL" />
            <COACH firstname="Jael" gender="F" lastname="Michel" />
            <COACH firstname="Annick" gender="F" lastname="Willemsen" nation="NED" license="25170" />
          </COACHES>
        </CLUB>
        <CLUB type="CLUB" code="STKP" nation="SUI" region="RZW" clubid="14172" name="Schwimmteam Kaiseraugst-Pratteln" name.en="Stkp" shortname="Stkp">
          <ATHLETES>
            <ATHLETE firstname="Lisa" lastname="Matter" birthdate="2011-01-02" gender="F" nation="SUI" athleteid="14183">
              <RESULTS>
                <RESULT eventid="1073" points="124" swimtime="00:00:51.28" resultid="14184" heatid="12875" lane="1" entrytime="00:00:54.00" />
                <RESULT eventid="1092" points="120" swimtime="00:00:57.83" resultid="14185" heatid="12888" lane="3" entrytime="00:01:02.00" />
                <RESULT eventid="1106" points="127" swimtime="00:00:45.55" resultid="14186" heatid="12916" lane="4" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olivia" lastname="Zurflueh" birthdate="2012-10-10" gender="F" nation="SUI" athleteid="14203">
              <RESULTS>
                <RESULT eventid="1073" points="133" swimtime="00:00:50.13" resultid="14204" heatid="12875" lane="3" entrytime="00:00:54.00" />
                <RESULT eventid="1092" points="128" swimtime="00:00:56.55" resultid="14205" heatid="12890" lane="2" entrytime="00:00:59.00" />
                <RESULT eventid="1106" points="129" swimtime="00:00:45.32" resultid="14206" heatid="12915" lane="3" entrytime="00:00:48.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Weichsel" birthdate="2010-08-31" gender="F" nation="SUI" athleteid="14199">
              <RESULTS>
                <RESULT eventid="1065" points="117" swimtime="00:01:51.97" resultid="14200" heatid="12859" lane="2" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="123" swimtime="00:02:05.26" resultid="14201" heatid="12898" lane="1" entrytime="00:01:59.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="121" swimtime="00:01:41.39" resultid="14202" heatid="12926" lane="2" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Thea" lastname="Richards" birthdate="2010-04-12" gender="F" nation="GBR" athleteid="14187">
              <RESULTS>
                <RESULT eventid="1065" points="125" swimtime="00:01:49.73" resultid="14188" heatid="12859" lane="1" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="127" swimtime="00:01:39.87" resultid="14189" heatid="12927" lane="4" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vangelis" lastname="Markopoulos" birthdate="2005-11-24" gender="M" nation="SUI" license="119737" athleteid="14178">
              <RESULTS>
                <RESULT eventid="1141" status="WDR" swimtime="00:00:00.00" resultid="14179" heatid="12973" lane="4" entrytime="00:01:28.00" />
                <RESULT eventid="1161" status="WDR" swimtime="00:00:00.00" resultid="14180" heatid="13004" lane="1" entrytime="00:02:50.00" />
                <RESULT eventid="1171" status="WDR" swimtime="00:00:00.00" resultid="14181" heatid="13014" lane="3" entrytime="00:01:40.00" />
                <RESULT eventid="1181" status="WDR" swimtime="00:00:00.00" resultid="14182" heatid="13035" lane="1" entrytime="00:01:18.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filip" lastname="Dokic" birthdate="2007-05-03" gender="M" nation="BIH" license="106113" athleteid="14173">
              <RESULTS>
                <RESULT eventid="1131" points="164" swimtime="00:01:27.28" resultid="14174" heatid="12957" lane="2" entrytime="00:01:26.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="223" swimtime="00:01:21.15" resultid="14175" heatid="12993" lane="3" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1161" points="251" swimtime="00:02:37.53" resultid="14176" heatid="13004" lane="2" entrytime="00:02:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.56" />
                    <SPLIT distance="100" swimtime="00:01:16.26" />
                    <SPLIT distance="150" swimtime="00:01:59.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="283" swimtime="00:01:08.41" resultid="14177" heatid="13036" lane="2" entrytime="00:01:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna Sol" lastname="Tüller" birthdate="2007-11-08" gender="F" nation="SUI" athleteid="14195">
              <RESULTS>
                <RESULT eventid="1136" points="138" swimtime="00:01:46.12" resultid="14196" heatid="12962" lane="3" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1166" points="133" swimtime="00:02:02.16" resultid="14197" heatid="13007" lane="2" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="159" swimtime="00:01:32.61" resultid="14198" heatid="13019" lane="3" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sriraam" lastname="Sivasundaran" birthdate="2007-01-23" gender="M" nation="SUI" license="110585" athleteid="14190">
              <RESULTS>
                <RESULT eventid="1141" points="153" swimtime="00:01:30.36" resultid="14191" heatid="12971" lane="3" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="170" swimtime="00:01:28.79" resultid="14192" heatid="12991" lane="4" entrytime="00:01:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1161" points="153" swimtime="00:03:05.72" resultid="14193" heatid="13003" lane="2" entrytime="00:02:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.59" />
                    <SPLIT distance="100" swimtime="00:01:25.36" />
                    <SPLIT distance="150" swimtime="00:02:15.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="152" swimtime="00:01:24.12" resultid="14194" heatid="13033" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SRSO" nation="SUI" region="RZW" clubid="11718" name="Swim Regio Solothurn">
          <ATHLETES>
            <ATHLETE firstname="Anna" lastname="Blazek" birthdate="2008-01-17" gender="F" nation="SUI" license="107521" athleteid="13640">
              <RESULTS>
                <RESULT eventid="1125" points="389" swimtime="00:01:14.77" resultid="13641" heatid="12953" lane="2" entrytime="00:01:15.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="403" swimtime="00:02:29.45" resultid="13642" heatid="12999" lane="1" entrytime="00:02:32.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.36" />
                    <SPLIT distance="100" swimtime="00:01:12.11" />
                    <SPLIT distance="150" swimtime="00:01:51.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="390" swimtime="00:01:08.74" resultid="13643" heatid="13024" lane="4" entrytime="00:01:10.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Levi" lastname="Berger" birthdate="2013-04-03" gender="M" nation="SUI" athleteid="13630">
              <RESULTS>
                <RESULT eventid="1076" points="41" swimtime="00:01:04.02" resultid="13631" heatid="12879" lane="1" entrytime="00:01:05.52" />
                <RESULT eventid="1109" points="34" swimtime="00:01:01.77" resultid="13632" heatid="12919" lane="2" entrytime="00:01:08.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alen" lastname="Besirovic" birthdate="2011-08-05" gender="M" nation="SUI" athleteid="13633">
              <RESULTS>
                <RESULT eventid="1076" points="51" swimtime="00:00:59.87" resultid="13634" heatid="12878" lane="2" entrytime="00:01:15.00" />
                <RESULT eventid="1109" points="53" swimtime="00:00:53.40" resultid="13635" heatid="12920" lane="4" entrytime="00:01:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Samuel" lastname="Kaiser" birthdate="2006-02-20" gender="M" nation="SUI" license="101209" athleteid="13694">
              <RESULTS>
                <RESULT eventid="1151" points="359" swimtime="00:01:09.28" resultid="13695" heatid="12995" lane="3" entrytime="00:01:17.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="410" swimtime="00:01:14.48" resultid="13696" heatid="13018" lane="3" entrytime="00:01:14.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caroline Mathilde" lastname="Bang" birthdate="2006-10-15" gender="F" nation="DEN" license="116476" athleteid="13628">
              <RESULTS>
                <RESULT eventid="1146" points="405" swimtime="00:01:16.33" resultid="13629" heatid="12990" lane="1" entrytime="00:01:10.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matej" lastname="Niznik" birthdate="2009-01-20" gender="M" nation="SVK" athleteid="13708">
              <RESULTS>
                <RESULT eventid="1070" points="133" swimtime="00:01:34.68" resultid="13709" heatid="12865" lane="2" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="201" swimtime="00:01:34.43" resultid="13710" heatid="12909" lane="4" entrytime="00:01:53.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="188" swimtime="00:01:18.38" resultid="13711" heatid="12938" lane="1" entrytime="00:01:40.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valentino" lastname="Tamburino" birthdate="2008-02-24" gender="M" nation="SUI" license="107843" athleteid="13727">
              <RESULTS>
                <RESULT eventid="1141" points="353" swimtime="00:01:08.38" resultid="13728" heatid="12977" lane="1" entrytime="00:01:09.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="330" swimtime="00:01:11.29" resultid="13729" heatid="12993" lane="2" entrytime="00:01:23.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="395" swimtime="00:01:01.20" resultid="13730" heatid="13040" lane="4" entrytime="00:01:01.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Noah" lastname="Schärer" birthdate="2007-01-30" gender="M" nation="SUI" license="122145" athleteid="13712">
              <RESULTS>
                <RESULT eventid="1151" points="385" swimtime="00:01:07.70" resultid="13713" heatid="12994" lane="1" entrytime="00:01:21.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="381" swimtime="00:01:16.33" resultid="13714" heatid="13015" lane="3" entrytime="00:01:30.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jana" lastname="Brunner" birthdate="2005-08-20" gender="F" nation="SUI" license="105642" athleteid="13644">
              <RESULTS>
                <RESULT eventid="1146" points="437" swimtime="00:01:14.42" resultid="13645" heatid="12989" lane="3" entrytime="00:01:14.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1166" points="395" swimtime="00:01:24.98" resultid="13646" heatid="14115" lane="4" entrytime="00:01:21.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="418" swimtime="00:01:07.16" resultid="13647" heatid="13030" lane="1" entrytime="00:01:04.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giada" lastname="Cuda" birthdate="2007-05-17" gender="F" nation="SUI" license="112149" athleteid="13668">
              <RESULTS>
                <RESULT eventid="1125" points="408" swimtime="00:01:13.57" resultid="13669" heatid="12954" lane="4" entrytime="00:01:15.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="432" swimtime="00:01:14.70" resultid="13670" heatid="12986" lane="2" entrytime="00:01:18.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1166" points="440" swimtime="00:01:21.95" resultid="13671" heatid="14115" lane="1" entrytime="00:01:21.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giulia Sarai" lastname="Günther" birthdate="2011-11-29" gender="F" nation="SUI" license="121779" athleteid="13672">
              <RESULTS>
                <RESULT eventid="1073" points="75" swimtime="00:01:00.64" resultid="13673" heatid="12871" lane="2" entrytime="00:01:15.00" />
                <RESULT eventid="1092" points="98" swimtime="00:01:01.87" resultid="13674" heatid="12886" lane="2" entrytime="00:01:20.00" />
                <RESULT eventid="1106" points="74" swimtime="00:00:54.55" resultid="13675" heatid="12912" lane="2" entrytime="00:01:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valerie Anna" lastname="Laeubli" birthdate="2010-03-03" gender="F" nation="SUI" license="120075" athleteid="13697">
              <RESULTS>
                <RESULT eventid="1065" points="218" swimtime="00:01:31.08" resultid="13698" heatid="12857" lane="1" entrytime="00:01:58.65" />
                <RESULT eventid="1099" points="217" swimtime="00:01:43.69" resultid="13699" heatid="12900" lane="1" entrytime="00:01:53.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="246" swimtime="00:01:20.19" resultid="13700" heatid="12926" lane="1" entrytime="00:01:49.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stefanie" lastname="Christen" birthdate="2009-01-30" gender="F" nation="SUI" license="107842" athleteid="13664">
              <RESULTS>
                <RESULT eventid="1099" points="324" swimtime="00:01:30.79" resultid="13665" heatid="12904" lane="2" entrytime="00:01:26.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1053" points="233" swimtime="00:00:39.61" resultid="13666" heatid="12849" lane="2" entrytime="00:00:41.66" entrycourse="LCM" />
                <RESULT eventid="1112" points="294" swimtime="00:01:15.52" resultid="13667" heatid="12934" lane="3" entrytime="00:01:13.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vania" lastname="von Känel" birthdate="2012-12-23" gender="F" nation="SUI" athleteid="13731">
              <RESULTS>
                <RESULT eventid="1073" points="109" swimtime="00:00:53.51" resultid="13732" heatid="12871" lane="3" entrytime="00:01:15.00" />
                <RESULT eventid="1106" points="85" swimtime="00:00:52.03" resultid="13733" heatid="12912" lane="3" entrytime="00:01:10.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mira" lastname="Leibundgut" birthdate="2008-09-20" gender="F" nation="SUI" license="107744" athleteid="13704">
              <RESULTS>
                <RESULT eventid="1125" points="326" swimtime="00:01:19.34" resultid="13705" heatid="12953" lane="4" entrytime="00:01:18.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="407" swimtime="00:02:28.91" resultid="13706" heatid="13000" lane="3" entrytime="00:02:25.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.66" />
                    <SPLIT distance="100" swimtime="00:01:12.66" />
                    <SPLIT distance="150" swimtime="00:01:51.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="387" swimtime="00:01:08.91" resultid="13707" heatid="13029" lane="4" entrytime="00:01:05.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Jost" birthdate="2005-04-19" gender="F" nation="SUI" license="37019" athleteid="13686">
              <RESULTS>
                <RESULT eventid="1125" points="445" swimtime="00:01:11.48" resultid="13687" heatid="12955" lane="4" entrytime="00:01:09.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="417" swimtime="00:01:15.59" resultid="13688" heatid="12989" lane="2" entrytime="00:01:13.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="424" swimtime="00:01:06.88" resultid="13689" heatid="13030" lane="4" entrytime="00:01:04.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dario" lastname="Burkhalter" birthdate="2009-10-29" gender="M" nation="SUI" athleteid="13652">
              <RESULTS>
                <RESULT eventid="1070" points="108" swimtime="00:01:41.19" resultid="13653" heatid="12867" lane="4" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="140" swimtime="00:01:46.36" resultid="13654" heatid="12909" lane="3" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="128" swimtime="00:01:29.17" resultid="13655" heatid="12938" lane="2" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Seraina" lastname="Häfliger" birthdate="2012-08-14" gender="F" nation="SUI" athleteid="13676">
              <RESULTS>
                <RESULT eventid="1073" points="116" swimtime="00:00:52.42" resultid="13677" heatid="12875" lane="4" entrytime="00:00:54.24" />
                <RESULT eventid="1106" points="101" swimtime="00:00:49.11" resultid="13678" heatid="12914" lane="3" entrytime="00:00:50.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Melanie" lastname="Christen" birthdate="2011-10-04" gender="F" nation="SUI" license="116469" athleteid="13660">
              <RESULTS>
                <RESULT eventid="1073" points="137" swimtime="00:00:49.65" resultid="13661" heatid="12872" lane="3" entrytime="00:01:00.00" />
                <RESULT eventid="1092" points="151" swimtime="00:00:53.54" resultid="13662" heatid="12887" lane="2" entrytime="00:01:06.09" />
                <RESULT eventid="1106" points="117" swimtime="00:00:46.83" resultid="13663" heatid="12913" lane="1" entrytime="00:00:57.19" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lea" lastname="Würgler" birthdate="2009-06-29" gender="F" nation="SUI" athleteid="13734">
              <RESULTS>
                <RESULT eventid="1065" points="127" swimtime="00:01:48.99" resultid="13735" heatid="12859" lane="3" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="201" swimtime="00:01:46.38" resultid="13736" heatid="12897" lane="4" entrytime="00:02:08.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="177" swimtime="00:01:29.37" resultid="13737" heatid="12927" lane="1" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eliott" lastname="André" birthdate="2007-10-13" gender="M" nation="SUI" athleteid="13624">
              <RESULTS>
                <RESULT eventid="1141" points="176" swimtime="00:01:26.14" resultid="13625" heatid="12972" lane="2" entrytime="00:01:30.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="165" swimtime="00:01:40.86" resultid="13626" heatid="13013" lane="3" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="223" swimtime="00:01:14.03" resultid="13627" heatid="13036" lane="1" entrytime="00:01:14.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valérie" lastname="Chiesa" birthdate="2007-02-21" gender="F" nation="SUI" license="113151" athleteid="13656">
              <RESULTS>
                <RESULT eventid="1146" points="342" swimtime="00:01:20.80" resultid="13657" heatid="12979" lane="3" entrytime="00:01:37.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1166" points="342" swimtime="00:01:29.09" resultid="13658" heatid="13011" lane="3" entrytime="00:01:29.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="349" swimtime="00:01:11.32" resultid="13659" heatid="13027" lane="2" entrytime="00:01:07.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tim" lastname="Honsberger" birthdate="2008-08-08" gender="M" nation="SUI" athleteid="13682">
              <RESULTS>
                <RESULT comment="209 - Zehen beider Füsse nicht in Kontakt mit Wand oder Anschlagplatte (Start)" eventid="1141" status="DSQ" swimtime="00:01:26.38" resultid="13683" heatid="12970" lane="2" entrytime="00:01:44.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="153" swimtime="00:01:43.41" resultid="13684" heatid="13013" lane="1" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="231" swimtime="00:01:13.14" resultid="13685" heatid="13034" lane="3" entrytime="00:01:18.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hannah" lastname="Kaiser" birthdate="2009-02-11" gender="F" nation="SUI" license="108993" athleteid="13690">
              <RESULTS>
                <RESULT eventid="1065" points="158" swimtime="00:01:41.50" resultid="13691" heatid="12861" lane="2" entrytime="00:01:38.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="189" swimtime="00:01:48.57" resultid="13692" heatid="12899" lane="1" entrytime="00:01:55.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="165" swimtime="00:01:31.47" resultid="13693" heatid="12928" lane="4" entrytime="00:01:38.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Xenia" lastname="Signoroni" birthdate="2005-11-16" gender="F" nation="SUI" license="37039" athleteid="13715">
              <RESULTS>
                <RESULT eventid="1125" points="371" swimtime="00:01:15.97" resultid="13716" heatid="12955" lane="1" entrytime="00:01:09.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="354" swimtime="00:01:17.53" resultid="13717" heatid="12968" lane="2" entrytime="00:01:11.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="412" swimtime="00:01:07.50" resultid="13718" heatid="13030" lane="2" entrytime="00:01:04.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lena" lastname="Leibundgut" birthdate="2004-08-26" gender="F" nation="SUI" license="36311" athleteid="13701">
              <RESULTS>
                <RESULT eventid="1125" points="489" swimtime="00:01:09.29" resultid="13702" heatid="12955" lane="2" entrytime="00:01:08.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="570" swimtime="00:02:13.14" resultid="13703" heatid="13001" lane="2" entrytime="00:02:09.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.60" />
                    <SPLIT distance="100" swimtime="00:01:05.16" />
                    <SPLIT distance="150" swimtime="00:01:39.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mailey Sue" lastname="Bruns" birthdate="2011-09-12" gender="F" nation="GER" license="120076" athleteid="13648">
              <RESULTS>
                <RESULT eventid="1073" points="242" swimtime="00:00:41.04" resultid="13649" heatid="12876" lane="3" entrytime="00:00:52.00" />
                <RESULT eventid="1092" points="174" swimtime="00:00:51.14" resultid="13650" heatid="12889" lane="1" entrytime="00:01:00.00" />
                <RESULT eventid="1106" points="251" swimtime="00:00:36.31" resultid="13651" heatid="12915" lane="2" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tobias" lastname="Birrer" birthdate="2008-05-21" gender="M" nation="SUI" license="107520" athleteid="13636">
              <RESULTS>
                <RESULT eventid="1131" points="278" swimtime="00:01:13.16" resultid="13637" heatid="12960" lane="2" entrytime="00:01:13.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="319" swimtime="00:01:12.05" resultid="13638" heatid="12994" lane="3" entrytime="00:01:21.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="293" swimtime="00:01:23.24" resultid="13639" heatid="13017" lane="1" entrytime="00:01:22.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tamara" lastname="Stooss" birthdate="2008-03-10" gender="F" nation="SUI" license="109133" athleteid="13719">
              <RESULTS>
                <RESULT eventid="1125" points="323" swimtime="00:01:19.52" resultid="13720" heatid="12953" lane="3" entrytime="00:01:16.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="377" swimtime="00:01:18.19" resultid="13721" heatid="12982" lane="2" entrytime="00:01:25.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="441" swimtime="00:01:06.01" resultid="13722" heatid="13029" lane="2" entrytime="00:01:04.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1122" points="82" swimtime="00:03:07.62" resultid="13738" heatid="12948" lane="1" entrytime="00:03:26.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.07" />
                    <SPLIT distance="100" swimtime="00:01:14.27" />
                    <SPLIT distance="150" swimtime="00:02:06.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13708" number="1" />
                    <RELAYPOSITION athleteid="13652" number="2" />
                    <RELAYPOSITION athleteid="13633" number="3" />
                    <RELAYPOSITION athleteid="13630" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1191" points="458" swimtime="00:03:57.37" resultid="13739" heatid="13045" lane="2" entrytime="00:04:02.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.71" />
                    <SPLIT distance="100" swimtime="00:01:00.09" />
                    <SPLIT distance="150" swimtime="00:01:29.45" />
                    <SPLIT distance="200" swimtime="00:02:01.46" />
                    <SPLIT distance="250" swimtime="00:02:29.71" />
                    <SPLIT distance="300" swimtime="00:03:01.79" />
                    <SPLIT distance="350" swimtime="00:03:28.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13694" number="1" />
                    <RELAYPOSITION athleteid="13636" number="2" />
                    <RELAYPOSITION athleteid="13727" number="3" />
                    <RELAYPOSITION athleteid="13712" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1119" points="250" swimtime="00:02:26.82" resultid="13740" heatid="12946" lane="3" entrytime="00:02:50.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                    <SPLIT distance="100" swimtime="00:01:14.27" />
                    <SPLIT distance="150" swimtime="00:01:53.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13697" number="1" />
                    <RELAYPOSITION athleteid="13734" number="2" />
                    <RELAYPOSITION athleteid="13690" number="3" />
                    <RELAYPOSITION athleteid="13664" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1186" points="521" swimtime="00:04:16.60" resultid="13741" heatid="13043" lane="3" entrytime="00:04:09.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.57" />
                    <SPLIT distance="100" swimtime="00:01:04.31" />
                    <SPLIT distance="150" swimtime="00:01:35.82" />
                    <SPLIT distance="200" swimtime="00:02:10.57" />
                    <SPLIT distance="250" swimtime="00:02:41.78" />
                    <SPLIT distance="300" swimtime="00:03:15.25" />
                    <SPLIT distance="350" swimtime="00:03:44.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13628" number="1" />
                    <RELAYPOSITION athleteid="13686" number="2" />
                    <RELAYPOSITION athleteid="13719" number="3" />
                    <RELAYPOSITION athleteid="13701" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1119" points="116" swimtime="00:03:09.16" resultid="13742" heatid="12945" lane="3" entrytime="00:03:45.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.55" />
                    <SPLIT distance="100" swimtime="00:01:24.54" />
                    <SPLIT distance="150" swimtime="00:02:16.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13648" number="1" />
                    <RELAYPOSITION athleteid="13660" number="2" />
                    <RELAYPOSITION athleteid="13676" number="3" />
                    <RELAYPOSITION athleteid="13672" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1186" points="454" swimtime="00:04:28.68" resultid="13743" heatid="13042" lane="2" entrytime="00:04:23.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.56" />
                    <SPLIT distance="100" swimtime="00:01:06.14" />
                    <SPLIT distance="150" swimtime="00:01:38.13" />
                    <SPLIT distance="200" swimtime="00:02:12.93" />
                    <SPLIT distance="250" swimtime="00:02:45.38" />
                    <SPLIT distance="300" swimtime="00:03:21.57" />
                    <SPLIT distance="350" swimtime="00:03:53.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13644" number="1" />
                    <RELAYPOSITION athleteid="13715" number="2" />
                    <RELAYPOSITION athleteid="13668" number="3" />
                    <RELAYPOSITION athleteid="13704" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SVB" nation="SUI" region="RZW" clubid="12648" name="Schwimmverein beider Basel" shortname="SV Basel">
          <ATHLETES>
            <ATHLETE firstname="Marah Anaïs" lastname="Becht" birthdate="2009-06-19" gender="F" nation="SUI" license="120382" athleteid="14536">
              <RESULTS>
                <RESULT eventid="1065" points="315" swimtime="00:01:20.59" resultid="14537" heatid="12863" lane="3" entrytime="00:01:19.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="392" swimtime="00:01:08.63" resultid="14538" heatid="12935" lane="1" entrytime="00:01:08.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Niederfeld" birthdate="2009-01-01" gender="M" nation="SUI" license="112793" athleteid="14610">
              <RESULTS>
                <RESULT comment="204 - Starten vor dem Startkommando" eventid="1060" status="DSQ" swimtime="00:00:41.67" resultid="14611" heatid="12855" lane="4" entrytime="00:00:43.21" entrycourse="LCM" />
                <RESULT eventid="1103" points="133" swimtime="00:01:48.18" resultid="14612" heatid="12907" lane="3" entrytime="00:02:00.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="160" swimtime="00:01:22.65" resultid="14613" heatid="12939" lane="3" entrytime="00:01:32.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robin" lastname="Marc" birthdate="2008-09-15" gender="M" nation="SUI" athleteid="14598">
              <RESULTS>
                <RESULT eventid="1141" points="163" swimtime="00:01:28.30" resultid="14599" heatid="12972" lane="3" entrytime="00:01:31.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="179" swimtime="00:01:27.36" resultid="14600" heatid="12991" lane="3" entrytime="00:01:36.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="193" swimtime="00:01:17.72" resultid="14601" heatid="13035" lane="3" entrytime="00:01:17.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ernesto" lastname="Calgua" birthdate="2008-01-01" gender="M" nation="SUI" athleteid="14551">
              <RESULTS>
                <RESULT eventid="1141" points="170" swimtime="00:01:27.11" resultid="14552" heatid="12971" lane="2" entrytime="00:01:37.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.58" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="404 - Nicht in Rückenlage angeschlagen (Ziel)" eventid="1151" status="DSQ" swimtime="00:01:30.90" resultid="14553" heatid="12991" lane="2" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="228" swimtime="00:01:13.48" resultid="14554" heatid="13036" lane="4" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Annika" lastname="Scharbert" birthdate="2009-10-11" gender="F" nation="SUI" license="112799" athleteid="14634">
              <RESULTS>
                <RESULT eventid="1053" points="224" swimtime="00:00:40.12" resultid="14635" heatid="12848" lane="1" entrytime="00:00:49.65" entrycourse="SCM" />
                <RESULT eventid="1099" points="247" swimtime="00:01:39.28" resultid="14636" heatid="12903" lane="1" entrytime="00:01:39.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="250" swimtime="00:01:19.76" resultid="14637" heatid="12931" lane="2" entrytime="00:01:22.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miriam" lastname="Colzani" birthdate="2009-12-26" gender="F" nation="ITA" athleteid="14555">
              <RESULTS>
                <RESULT eventid="1053" points="235" swimtime="00:00:39.48" resultid="14556" heatid="12849" lane="1" entrytime="00:00:45.49" entrycourse="LCM" />
                <RESULT eventid="1099" points="229" swimtime="00:01:41.83" resultid="14557" heatid="12900" lane="4" entrytime="00:01:53.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="246" swimtime="00:01:20.11" resultid="14558" heatid="12931" lane="3" entrytime="00:01:23.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carl-Leopold" lastname="Hackner" birthdate="2010-02-26" gender="M" nation="SUI" athleteid="14570">
              <RESULTS>
                <RESULT eventid="1070" points="218" swimtime="00:01:20.25" resultid="14571" heatid="12868" lane="3" entrytime="00:01:24.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="187" swimtime="00:01:36.71" resultid="14572" heatid="12909" lane="1" entrytime="00:01:50.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="235" swimtime="00:01:12.76" resultid="14573" heatid="12942" lane="1" entrytime="00:01:14.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcos" lastname="Rivero" birthdate="2005-03-30" gender="M" nation="FRA" license="115177" athleteid="14630">
              <RESULTS>
                <RESULT eventid="1131" points="289" swimtime="00:01:12.20" resultid="14631" heatid="12958" lane="3" entrytime="00:01:21.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1161" points="368" swimtime="00:02:18.60" resultid="14632" heatid="13006" lane="1" entrytime="00:02:21.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.83" />
                    <SPLIT distance="100" swimtime="00:01:06.25" />
                    <SPLIT distance="150" swimtime="00:01:43.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="390" swimtime="00:01:01.48" resultid="14633" heatid="13039" lane="1" entrytime="00:01:03.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martha" lastname="Bolten" birthdate="2007-01-15" gender="F" nation="SUI" license="117350" athleteid="14543">
              <RESULTS>
                <RESULT eventid="1136" points="302" swimtime="00:01:21.75" resultid="14544" heatid="12965" lane="3" entrytime="00:01:26.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="354" swimtime="00:01:19.85" resultid="14545" heatid="12985" lane="4" entrytime="00:01:22.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="401" swimtime="00:01:08.13" resultid="14546" heatid="13026" lane="2" entrytime="00:01:07.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nina" lastname="Zangger" birthdate="2005-12-09" gender="F" nation="SUI" license="113156" athleteid="14646">
              <RESULTS>
                <RESULT eventid="1125" points="292" swimtime="00:01:22.29" resultid="14647" heatid="12950" lane="3" entrytime="00:01:29.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="358" swimtime="00:01:19.57" resultid="14648" heatid="12985" lane="1" entrytime="00:01:22.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="351" swimtime="00:01:11.21" resultid="14649" heatid="13024" lane="3" entrytime="00:01:10.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hector" lastname="Rivero" birthdate="2007-01-01" gender="M" nation="FRA" license="119209" athleteid="14626">
              <RESULTS>
                <RESULT eventid="1161" points="289" swimtime="00:02:30.17" resultid="14627" heatid="13005" lane="3" entrytime="00:02:27.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                    <SPLIT distance="100" swimtime="00:01:12.96" />
                    <SPLIT distance="150" swimtime="00:01:52.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="261" swimtime="00:01:10.24" resultid="14628" heatid="13037" lane="1" entrytime="00:01:07.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="200" swimtime="00:01:22.55" resultid="14629" heatid="12974" lane="4" entrytime="00:01:21.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laila Brooke" lastname="Niederfeld" birthdate="2007-02-15" gender="F" nation="GER" license="105814" athleteid="14606">
              <RESULTS>
                <RESULT eventid="1125" points="351" swimtime="00:01:17.35" resultid="14607" heatid="12953" lane="1" entrytime="00:01:17.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="361" swimtime="00:01:19.33" resultid="14608" heatid="12986" lane="4" entrytime="00:01:20.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="397" swimtime="00:01:08.37" resultid="14609" heatid="13026" lane="3" entrytime="00:01:08.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ella" lastname="Aebi" birthdate="2009-07-16" gender="F" nation="SUI" license="115169" athleteid="14520">
              <RESULTS>
                <RESULT eventid="1053" points="301" swimtime="00:00:36.35" resultid="14521" heatid="12850" lane="1" entrytime="00:00:41.09" entrycourse="LCM" />
                <RESULT eventid="1099" points="333" swimtime="00:01:29.92" resultid="14522" heatid="12904" lane="3" entrytime="00:01:29.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="366" swimtime="00:01:10.21" resultid="14523" heatid="12935" lane="4" entrytime="00:01:10.71" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Blake" lastname="Harada" birthdate="2008-04-05" gender="M" nation="SUI" license="119173" athleteid="14578">
              <RESULTS>
                <RESULT eventid="1131" points="177" swimtime="00:01:24.94" resultid="14579" heatid="12957" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="256" swimtime="00:01:17.60" resultid="14580" heatid="12992" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="242" swimtime="00:01:12.10" resultid="14581" heatid="13034" lane="2" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Duygu Naz" lastname="Aykut" birthdate="2008-02-04" gender="F" nation="SUI" license="116161" athleteid="14524">
              <RESULTS>
                <RESULT eventid="1136" points="302" swimtime="00:01:21.73" resultid="14525" heatid="12966" lane="1" entrytime="00:01:21.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="302" swimtime="00:01:24.19" resultid="14526" heatid="12980" lane="2" entrytime="00:01:31.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="328" swimtime="00:01:12.79" resultid="14527" heatid="13023" lane="1" entrytime="00:01:12.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Procopio" birthdate="2007-12-05" gender="F" nation="SUI" license="119121" athleteid="14618">
              <RESULTS>
                <RESULT eventid="1125" points="220" swimtime="00:01:30.45" resultid="14619" heatid="12950" lane="2" entrytime="00:01:28.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="274" swimtime="00:01:26.98" resultid="14620" heatid="12982" lane="3" entrytime="00:01:26.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="296" swimtime="00:01:15.32" resultid="14621" heatid="13022" lane="3" entrytime="00:01:14.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ann-Sophie" lastname="Baur" birthdate="2009-04-09" gender="F" nation="SUI" license="112734" athleteid="14532">
              <RESULTS>
                <RESULT eventid="1053" points="297" swimtime="00:00:36.52" resultid="14533" heatid="12851" lane="3" entrytime="00:00:38.74" entrycourse="LCM" />
                <RESULT eventid="1099" points="309" swimtime="00:01:32.24" resultid="14534" heatid="12904" lane="1" entrytime="00:01:33.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="321" swimtime="00:01:13.38" resultid="14535" heatid="12933" lane="2" entrytime="00:01:15.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giuliana" lastname="Gamboni" birthdate="2009-07-07" gender="F" nation="SUI" license="6400" athleteid="14563">
              <RESULTS>
                <RESULT eventid="1099" points="225" swimtime="00:01:42.42" resultid="14564" heatid="12901" lane="1" entrytime="00:01:48.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="179" swimtime="00:01:29.14" resultid="14565" heatid="12931" lane="4" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lilja" lastname="Hausmann" birthdate="2010-04-01" gender="F" nation="SUI" athleteid="14582">
              <RESULTS>
                <RESULT eventid="1065" points="189" swimtime="00:01:35.61" resultid="14583" heatid="12860" lane="4" entrytime="00:01:46.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="262" swimtime="00:01:37.36" resultid="14584" heatid="12903" lane="2" entrytime="00:01:38.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="204" swimtime="00:01:25.23" resultid="14585" heatid="12929" lane="2" entrytime="00:01:27.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Chiara" lastname="Kesselgruber" birthdate="2010-01-10" gender="F" nation="SUI" license="119162" athleteid="14590">
              <RESULTS>
                <RESULT eventid="1065" points="240" swimtime="00:01:28.25" resultid="14591" heatid="12862" lane="2" entrytime="00:01:33.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="223" swimtime="00:01:42.77" resultid="14592" heatid="12902" lane="4" entrytime="00:01:46.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="245" swimtime="00:01:20.24" resultid="14593" heatid="12930" lane="2" entrytime="00:01:24.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yann" lastname="Giorgetti" birthdate="2007-01-01" gender="M" nation="FRA" license="119729" athleteid="14566">
              <RESULTS>
                <RESULT eventid="1141" points="332" swimtime="00:01:09.79" resultid="14567" heatid="12977" lane="4" entrytime="00:01:11.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="308" swimtime="00:01:12.93" resultid="14568" heatid="12993" lane="1" entrytime="00:01:25.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="363" swimtime="00:01:02.95" resultid="14569" heatid="13039" lane="3" entrytime="00:01:03.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dusan" lastname="Radivojevic" birthdate="2007-09-18" gender="M" nation="SUI" license="109817" athleteid="14622">
              <RESULTS>
                <RESULT eventid="1141" status="WDR" swimtime="00:00:00.00" resultid="14623" entrytime="00:01:16.67" entrycourse="LCM" />
                <RESULT eventid="1151" status="WDR" swimtime="00:00:00.00" resultid="14624" entrytime="00:01:29.36" entrycourse="SCM" />
                <RESULT eventid="1171" status="WDR" swimtime="00:00:00.00" resultid="14625" entrytime="00:01:26.50" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anastasia" lastname="Hak" birthdate="2010-01-01" gender="F" nation="SUI" athleteid="14574">
              <RESULTS>
                <RESULT eventid="1065" points="403" swimtime="00:01:14.28" resultid="14575" heatid="12863" lane="2" entrytime="00:01:14.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="340" swimtime="00:01:29.32" resultid="14576" heatid="12900" lane="3" entrytime="00:01:52.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="419" swimtime="00:01:07.12" resultid="14577" heatid="12935" lane="3" entrytime="00:01:07.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patricia" lastname="Luther" birthdate="2007-01-01" gender="F" nation="SUI" athleteid="14594">
              <RESULTS>
                <RESULT eventid="1125" points="215" swimtime="00:01:31.13" resultid="14595" heatid="12949" lane="2" entrytime="00:01:32.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="325" swimtime="00:01:22.19" resultid="14596" heatid="12985" lane="3" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="396" swimtime="00:01:08.41" resultid="14597" heatid="13026" lane="1" entrytime="00:01:08.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kevin" lastname="Barron" birthdate="2009-12-02" gender="M" nation="SUI" athleteid="14528">
              <RESULTS>
                <RESULT comment="304 - Schwimmen in Bauchlage vor der Wende (Wende ...)" eventid="1070" status="DSQ" swimtime="00:01:39.26" resultid="14529" heatid="12867" lane="2" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="146" swimtime="00:01:45.00" resultid="14530" heatid="12909" lane="2" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="107" swimtime="00:01:34.60" resultid="14531" heatid="12940" lane="3" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mareen" lastname="Scharbert" birthdate="2009-10-11" gender="F" nation="SUI" license="112800" athleteid="14638">
              <RESULTS>
                <RESULT eventid="1065" points="164" swimtime="00:01:40.08" resultid="14639" heatid="12858" lane="3" entrytime="00:01:51.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="237" swimtime="00:01:40.74" resultid="14640" heatid="12901" lane="2" entrytime="00:01:47.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="159" swimtime="00:01:32.71" resultid="14641" heatid="12928" lane="1" entrytime="00:01:36.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nils" lastname="Borer" birthdate="2009-08-08" gender="M" nation="SUI" license="117624" athleteid="14547">
              <RESULTS>
                <RESULT eventid="1060" points="195" swimtime="00:00:37.48" resultid="14548" heatid="12855" lane="1" entrytime="00:00:41.37" entrycourse="LCM" />
                <RESULT eventid="1103" points="286" swimtime="00:01:23.93" resultid="14549" heatid="12910" lane="2" entrytime="00:01:25.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="261" swimtime="00:01:10.24" resultid="14550" heatid="12942" lane="2" entrytime="00:01:09.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jasmine" lastname="Hoog" birthdate="2007-03-18" gender="F" nation="SUI" license="102616" athleteid="14586">
              <RESULTS>
                <RESULT eventid="1125" points="389" swimtime="00:01:14.75" resultid="14587" heatid="12952" lane="2" entrytime="00:01:18.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="357" swimtime="00:01:19.60" resultid="14588" heatid="12984" lane="3" entrytime="00:01:23.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="379" swimtime="00:01:09.42" resultid="14589" heatid="13027" lane="3" entrytime="00:01:07.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juliette" lastname="Frederiksen" birthdate="2008-08-17" gender="F" nation="SUI" athleteid="14559">
              <RESULTS>
                <RESULT eventid="1136" points="230" swimtime="00:01:29.51" resultid="14560" heatid="12963" lane="2" entrytime="00:01:36.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="246" swimtime="00:01:30.12" resultid="14561" heatid="12978" lane="4" entrytime="00:01:48.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="238" swimtime="00:01:21.07" resultid="14562" heatid="13019" lane="1" entrytime="00:01:40.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lauren" lastname="Milnes" birthdate="2007-01-01" gender="F" nation="SUI" license="119165" athleteid="14602">
              <RESULTS>
                <RESULT eventid="1125" points="316" swimtime="00:01:20.12" resultid="14603" heatid="12952" lane="4" entrytime="00:01:21.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="375" swimtime="00:01:18.30" resultid="14604" heatid="12983" lane="2" entrytime="00:01:24.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="399" swimtime="00:01:08.24" resultid="14605" heatid="13028" lane="4" entrytime="00:01:07.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ghanima" lastname="Bekhit" birthdate="2008-04-22" gender="F" nation="SUI" license="112795" athleteid="14539">
              <RESULTS>
                <RESULT eventid="1125" points="301" swimtime="00:01:21.45" resultid="14540" heatid="12951" lane="4" entrytime="00:01:27.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.34" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="204 - Starten vor dem Startkommando" eventid="1146" status="DSQ" swimtime="00:01:21.45" resultid="14541" heatid="12981" lane="1" entrytime="00:01:29.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="312" swimtime="00:01:14.07" resultid="14542" heatid="13024" lane="1" entrytime="00:01:10.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Palombi" birthdate="2009-02-12" gender="F" nation="ITA" athleteid="14614">
              <RESULTS>
                <RESULT eventid="1065" points="182" swimtime="00:01:36.72" resultid="14615" heatid="12860" lane="3" entrytime="00:01:43.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="217" swimtime="00:01:43.70" resultid="14616" heatid="12901" lane="4" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="228" swimtime="00:01:22.24" resultid="14617" heatid="12931" lane="1" entrytime="00:01:23.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cynthia" lastname="Wiedemann" birthdate="2005-09-19" gender="F" nation="SUI" license="7599" athleteid="14642">
              <RESULTS>
                <RESULT eventid="1146" points="383" swimtime="00:01:17.80" resultid="14643" heatid="12984" lane="2" entrytime="00:01:22.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="400" swimtime="00:02:29.80" resultid="14644" heatid="13000" lane="4" entrytime="00:02:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.65" />
                    <SPLIT distance="100" swimtime="00:01:11.59" />
                    <SPLIT distance="150" swimtime="00:01:51.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="418" swimtime="00:01:07.17" resultid="14645" heatid="13028" lane="1" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1122" points="196" swimtime="00:02:20.70" resultid="14650" heatid="14668" lane="2" entrytime="00:02:19.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.15" />
                    <SPLIT distance="100" swimtime="00:01:09.55" />
                    <SPLIT distance="150" swimtime="00:01:49.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14570" number="1" />
                    <RELAYPOSITION athleteid="14610" number="2" />
                    <RELAYPOSITION athleteid="14528" number="3" />
                    <RELAYPOSITION athleteid="14547" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1119" points="393" swimtime="00:02:06.27" resultid="14651" heatid="14669" lane="3" entrytime="00:02:14.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.91" />
                    <SPLIT distance="100" swimtime="00:01:05.42" />
                    <SPLIT distance="150" swimtime="00:01:36.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14536" number="1" />
                    <RELAYPOSITION athleteid="14532" number="2" />
                    <RELAYPOSITION athleteid="14520" number="3" />
                    <RELAYPOSITION athleteid="14574" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1119" points="256" swimtime="00:02:25.61" resultid="14652" heatid="14669" lane="4" entrytime="00:02:26.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.70" />
                    <SPLIT distance="100" swimtime="00:01:11.56" />
                    <SPLIT distance="150" swimtime="00:01:49.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14555" number="1" />
                    <RELAYPOSITION athleteid="14590" number="2" />
                    <RELAYPOSITION athleteid="14563" number="3" />
                    <RELAYPOSITION athleteid="14614" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SBO" nation="SUI" region="RZW" clubid="12336" name="Schwimmclub Bottmingen-Oberwil">
          <ATHLETES>
            <ATHLETE firstname="Magnus" lastname="Klein" birthdate="2011-05-02" gender="M" nation="SUI" athleteid="12384">
              <RESULTS>
                <RESULT eventid="1060" points="84" swimtime="00:00:49.63" resultid="12385" heatid="12853" lane="2" entrytime="00:00:51.90" />
                <RESULT eventid="1096" points="99" swimtime="00:00:54.54" resultid="12386" heatid="12895" lane="3" entrytime="00:00:51.49" />
                <RESULT comment="204 - Starten vor dem Startkommando" eventid="1109" status="DSQ" swimtime="00:00:39.50" resultid="12387" heatid="12923" lane="2" entrytime="00:00:40.02" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lena" lastname="Bur" birthdate="2012-05-01" gender="F" nation="SUI" athleteid="12359">
              <RESULTS>
                <RESULT eventid="1073" points="134" swimtime="00:00:49.96" resultid="12360" heatid="12877" lane="4" entrytime="00:00:50.77" />
                <RESULT eventid="1092" points="123" swimtime="00:00:57.30" resultid="12361" heatid="12891" lane="4" entrytime="00:00:58.82" />
                <RESULT eventid="1106" points="153" swimtime="00:00:42.80" resultid="12362" heatid="12914" lane="2" entrytime="00:00:49.29" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mark" lastname="Xu" birthdate="2009-09-01" gender="M" nation="GBR" athleteid="12449">
              <RESULTS>
                <RESULT eventid="1060" points="200" swimtime="00:00:37.15" resultid="12450" heatid="12855" lane="3" entrytime="00:00:41.02" />
                <RESULT eventid="1088" points="203" swimtime="00:02:48.97" resultid="12451" heatid="12884" lane="2" entrytime="00:03:00.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.34" />
                    <SPLIT distance="100" swimtime="00:01:18.38" />
                    <SPLIT distance="150" swimtime="00:02:04.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="220" swimtime="00:01:14.37" resultid="12452" heatid="12942" lane="4" entrytime="00:01:18.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henry" lastname="Von Girsewald" birthdate="2011-09-17" gender="M" nation="SUI" athleteid="12444">
              <RESULTS>
                <RESULT comment="204 - Starten vor dem Startkommando" eventid="1060" status="DSQ" swimtime="00:00:45.52" resultid="12445" heatid="12853" lane="3" entrytime="00:00:53.90" />
                <RESULT eventid="1076" points="110" swimtime="00:00:46.24" resultid="12446" heatid="12881" lane="3" entrytime="00:00:56.59" />
                <RESULT eventid="1096" points="103" swimtime="00:00:53.73" resultid="12447" heatid="12895" lane="4" entrytime="00:00:54.58" />
                <RESULT eventid="1109" points="123" swimtime="00:00:40.49" resultid="12448" heatid="12923" lane="4" entrytime="00:00:41.67" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jonathan" lastname="Ng" birthdate="2010-02-18" gender="M" nation="CAN" athleteid="12412">
              <RESULTS>
                <RESULT eventid="1070" status="WDR" swimtime="00:00:00.00" resultid="12413" heatid="12864" lane="1" />
                <RESULT eventid="1103" status="WDR" swimtime="00:00:00.00" resultid="12414" heatid="12906" lane="1" />
                <RESULT eventid="1116" status="WDR" swimtime="00:00:00.00" resultid="12415" heatid="12937" lane="4" entrytime="00:01:48.98" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Batu" lastname="Yüksel" birthdate="2013-12-25" gender="M" nation="TUR" athleteid="12453">
              <RESULTS>
                <RESULT eventid="1076" points="54" swimtime="00:00:58.47" resultid="12454" heatid="12878" lane="1" />
                <RESULT comment="403 - Nicht mit beiden Händen gleichzeitig angeschlagen (Ziel)" eventid="1096" status="DSQ" swimtime="00:01:23.12" resultid="12455" heatid="12892" lane="4" />
                <RESULT eventid="1109" points="40" swimtime="00:00:58.56" resultid="12456" heatid="12919" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elias" lastname="Mussio" birthdate="2004-11-04" gender="M" nation="SUI" license="46917" athleteid="12408">
              <RESULTS>
                <RESULT eventid="1171" points="423" swimtime="00:01:13.72" resultid="12409" heatid="13018" lane="1" entrytime="00:01:15.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="368" swimtime="00:01:06.66" resultid="12410" heatid="14653" lane="1" entrytime="00:01:07.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="434" swimtime="00:01:05.08" resultid="12411" heatid="12997" lane="1" entrytime="00:01:08.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tobi" lastname="Schnyder" birthdate="2007-07-05" gender="M" nation="SUI" athleteid="12420">
              <RESULTS>
                <RESULT eventid="1151" points="194" swimtime="00:01:25.06" resultid="12421" heatid="12992" lane="1" entrytime="00:01:30.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="217" swimtime="00:01:31.96" resultid="12422" heatid="13014" lane="2" entrytime="00:01:36.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="223" swimtime="00:01:14.02" resultid="12423" heatid="13035" lane="2" entrytime="00:01:16.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milla" lastname="Spielmann" birthdate="2008-07-19" gender="F" nation="SUI" license="110216" athleteid="12428">
              <RESULTS>
                <RESULT eventid="1136" points="297" swimtime="00:01:22.24" resultid="12429" heatid="12965" lane="2" entrytime="00:01:25.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="296" swimtime="00:02:45.62" resultid="12430" heatid="12998" lane="3" entrytime="00:03:12.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.46" />
                    <SPLIT distance="100" swimtime="00:01:19.92" />
                    <SPLIT distance="150" swimtime="00:02:03.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="280" swimtime="00:01:16.76" resultid="12431" heatid="13020" lane="2" entrytime="00:01:20.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Len" lastname="Goeppert" birthdate="2002-11-07" gender="M" nation="SUI" license="29782" athleteid="12371">
              <RESULTS>
                <RESULT eventid="1141" points="399" swimtime="00:01:05.61" resultid="12372" heatid="12970" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1161" points="463" swimtime="00:02:08.42" resultid="12373" heatid="13003" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.72" />
                    <SPLIT distance="100" swimtime="00:01:02.28" />
                    <SPLIT distance="150" swimtime="00:01:35.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="498" swimtime="00:00:56.69" resultid="12374" heatid="13033" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mathilde" lastname="Fredersdorf" birthdate="2008-05-26" gender="F" nation="SUI" license="110210" athleteid="12367">
              <RESULTS>
                <RESULT eventid="1125" points="372" swimtime="00:01:15.90" resultid="12368" heatid="12950" lane="4" entrytime="00:01:30.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="441" swimtime="00:01:14.19" resultid="12369" heatid="12983" lane="3" entrytime="00:01:24.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1166" points="416" swimtime="00:01:23.47" resultid="12370" heatid="13010" lane="3" entrytime="00:01:31.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Soufian" lastname="Beltman" birthdate="2009-04-28" gender="M" nation="NED" athleteid="12350">
              <RESULTS>
                <RESULT eventid="1060" points="109" swimtime="00:00:45.53" resultid="12351" heatid="12854" lane="1" entrytime="00:00:45.24" />
                <RESULT eventid="1088" points="142" swimtime="00:03:10.18" resultid="12352" heatid="12884" lane="4" entrytime="00:03:10.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.30" />
                    <SPLIT distance="100" swimtime="00:01:30.33" />
                    <SPLIT distance="150" swimtime="00:02:21.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="141" swimtime="00:01:26.24" resultid="12353" heatid="12941" lane="4" entrytime="00:01:24.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Florian" lastname="Barthlott" birthdate="2002-09-06" gender="M" nation="SUI" license="113867" athleteid="12337">
              <RESULTS>
                <RESULT eventid="1141" points="277" swimtime="00:01:14.11" resultid="12338" heatid="12975" lane="2" entrytime="00:01:13.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1161" points="383" swimtime="00:02:16.81" resultid="12339" heatid="13006" lane="3" entrytime="00:02:18.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.76" />
                    <SPLIT distance="100" swimtime="00:01:04.81" />
                    <SPLIT distance="150" swimtime="00:01:40.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="391" swimtime="00:01:01.41" resultid="12340" heatid="13039" lane="2" entrytime="00:01:02.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felix" lastname="Bayer" birthdate="2010-02-08" gender="M" nation="SUI" athleteid="12346">
              <RESULTS>
                <RESULT eventid="1070" points="144" swimtime="00:01:32.19" resultid="12347" heatid="12866" lane="4" entrytime="00:01:44.86" />
                <RESULT eventid="1103" points="154" swimtime="00:01:43.22" resultid="12348" heatid="12910" lane="1" entrytime="00:01:45.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="190" swimtime="00:01:18.11" resultid="12349" heatid="12941" lane="1" entrytime="00:01:20.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luc" lastname="Montavon" birthdate="2010-05-29" gender="M" nation="SUI" athleteid="12404">
              <RESULTS>
                <RESULT eventid="1070" points="66" swimtime="00:01:59.33" resultid="12405" heatid="12865" lane="4" entrytime="00:02:04.81">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.56" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="303 - Nicht mit beiden Händen gleichzeitig angeschlagen (Wende  ...)" eventid="1103" status="DSQ" swimtime="00:02:02.58" resultid="12406" heatid="12907" lane="1" entrytime="00:02:00.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="91" swimtime="00:01:39.72" resultid="12407" heatid="12937" lane="1" entrytime="00:01:45.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emma Sophie" lastname="Bayer" birthdate="2012-01-06" gender="F" nation="DEN" athleteid="12341">
              <RESULTS>
                <RESULT eventid="1053" points="113" swimtime="00:00:50.33" resultid="12342" heatid="12847" lane="3" entrytime="00:00:52.02" />
                <RESULT eventid="1073" points="108" swimtime="00:00:53.68" resultid="12343" heatid="12876" lane="2" entrytime="00:00:50.82" />
                <RESULT eventid="1092" points="210" swimtime="00:00:47.98" resultid="12344" heatid="14113" lane="2" entrytime="00:00:51.45" />
                <RESULT eventid="1106" points="181" swimtime="00:00:40.49" resultid="12345" heatid="12918" lane="2" entrytime="00:00:38.26" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Beltman" birthdate="2009-04-28" gender="F" nation="NED" athleteid="12354">
              <RESULTS>
                <RESULT eventid="1053" points="134" swimtime="00:00:47.62" resultid="12355" heatid="12848" lane="3" entrytime="00:00:48.27" />
                <RESULT eventid="1065" points="115" swimtime="00:01:52.79" resultid="12356" heatid="12858" lane="1" entrytime="00:01:53.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.88" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="206 - Unterwasserphase: Mehr als ein Delphinbeinschlag (Start)" eventid="1099" status="DSQ" swimtime="00:01:54.46" resultid="12357" heatid="12898" lane="4" entrytime="00:01:59.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="151" swimtime="00:01:34.30" resultid="12358" heatid="12935" lane="2" entrytime="00:00:31.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ruwen" lastname="Gu" birthdate="2010-04-28" gender="M" nation="CHN" athleteid="12379">
              <RESULTS>
                <RESULT eventid="1060" points="118" swimtime="00:00:44.22" resultid="12380" heatid="12853" lane="1" entrytime="00:00:54.02" />
                <RESULT eventid="1070" points="105" swimtime="00:01:42.22" resultid="12381" heatid="12866" lane="3" entrytime="00:01:42.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="135" swimtime="00:01:47.64" resultid="12382" heatid="12908" lane="3" entrytime="00:01:54.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="141" swimtime="00:01:26.30" resultid="12383" heatid="12939" lane="2" entrytime="00:01:30.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Linley" lastname="Mead" birthdate="2009-10-06" gender="F" nation="USA" athleteid="12400">
              <RESULTS>
                <RESULT eventid="1065" points="126" swimtime="00:01:49.22" resultid="12401" heatid="12859" lane="4" entrytime="00:01:50.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="139" swimtime="00:02:00.28" resultid="12402" heatid="12899" lane="3" entrytime="00:01:54.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="178" swimtime="00:01:29.25" resultid="12403" heatid="12929" lane="4" entrytime="00:01:28.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Moritz" lastname="Takes" birthdate="2010-01-01" gender="M" nation="GER" athleteid="12440">
              <RESULTS>
                <RESULT eventid="1060" points="119" swimtime="00:00:44.17" resultid="12441" heatid="12854" lane="2" entrytime="00:00:44.02" />
                <RESULT eventid="1070" points="155" swimtime="00:01:29.83" resultid="12442" heatid="12868" lane="4" entrytime="00:01:34.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="182" swimtime="00:01:19.25" resultid="12443" heatid="12941" lane="3" entrytime="00:01:20.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlotta" lastname="Diddoro" birthdate="2009-01-26" gender="F" nation="ITA" athleteid="12363">
              <RESULTS>
                <RESULT eventid="1065" points="110" swimtime="00:01:54.46" resultid="12364" heatid="12856" lane="2" entrytime="00:01:58.88" />
                <RESULT eventid="1099" points="162" swimtime="00:01:54.32" resultid="12365" heatid="12898" lane="3" entrytime="00:01:58.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="88" swimtime="00:01:52.76" resultid="12366" heatid="12925" lane="2" entrytime="00:01:52.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ruth" lastname="Leibfritz" birthdate="2012-01-17" gender="F" nation="GER" athleteid="12388">
              <RESULTS>
                <RESULT eventid="1073" points="88" swimtime="00:00:57.38" resultid="12389" heatid="12872" lane="1" entrytime="00:01:00.02" />
                <RESULT eventid="1092" points="106" swimtime="00:01:00.22" resultid="12390" heatid="12888" lane="1" entrytime="00:01:02.02" />
                <RESULT eventid="1106" points="104" swimtime="00:00:48.64" resultid="12391" heatid="12916" lane="1" entrytime="00:00:47.87" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Clara" lastname="Schwöbel" birthdate="2008-09-07" gender="F" nation="SUI" license="110220" athleteid="12424">
              <RESULTS>
                <RESULT eventid="1136" points="147" swimtime="00:01:43.92" resultid="12425" heatid="12963" lane="3" entrytime="00:01:42.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="178" swimtime="00:01:40.28" resultid="12426" heatid="12978" lane="2" entrytime="00:01:40.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1166" points="243" swimtime="00:01:39.88" resultid="12427" heatid="13008" lane="3" entrytime="00:01:45.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caspar" lastname="Takes" birthdate="2011-09-12" gender="M" nation="GER" athleteid="12436">
              <RESULTS>
                <RESULT eventid="1076" points="99" swimtime="00:00:47.90" resultid="12437" heatid="12882" lane="1" entrytime="00:00:50.46" />
                <RESULT eventid="1096" points="112" swimtime="00:00:52.32" resultid="12438" heatid="12895" lane="2" entrytime="00:00:51.48" />
                <RESULT eventid="1109" points="133" swimtime="00:00:39.49" resultid="12439" heatid="12923" lane="3" entrytime="00:00:40.02" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Oliver" lastname="Story" birthdate="2007-07-03" gender="M" nation="SUI" athleteid="12432">
              <RESULTS>
                <RESULT eventid="1141" points="163" swimtime="00:01:28.33" resultid="12433" heatid="12972" lane="1" entrytime="00:01:35.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1161" points="188" swimtime="00:02:53.43" resultid="12434" heatid="13003" lane="3" entrytime="00:02:55.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.38" />
                    <SPLIT distance="100" swimtime="00:01:20.77" />
                    <SPLIT distance="150" swimtime="00:02:07.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="197" swimtime="00:01:17.11" resultid="12435" heatid="13034" lane="1" entrytime="00:01:19.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lea" lastname="Gramke" birthdate="2006-07-04" gender="F" nation="SUI" license="110205" athleteid="12375">
              <RESULTS>
                <RESULT eventid="1136" points="483" swimtime="00:01:09.94" resultid="12376" heatid="12969" lane="1" entrytime="00:01:10.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="447" swimtime="00:01:11.42" resultid="12377" heatid="12954" lane="2" entrytime="00:01:10.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="477" swimtime="00:01:04.29" resultid="12378" heatid="13028" lane="2" entrytime="00:01:06.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1122" points="177" swimtime="00:02:25.42" resultid="12457" heatid="14668" lane="3" entrytime="00:02:30.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.31" />
                    <SPLIT distance="100" swimtime="00:01:13.46" />
                    <SPLIT distance="150" swimtime="00:01:49.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12346" number="1" />
                    <RELAYPOSITION athleteid="12379" number="2" />
                    <RELAYPOSITION athleteid="12440" number="3" />
                    <RELAYPOSITION athleteid="12350" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1191" points="400" swimtime="00:04:08.40" resultid="12458" heatid="13044" lane="2" entrytime="00:04:13.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.89" />
                    <SPLIT distance="100" swimtime="00:00:57.91" />
                    <SPLIT distance="150" swimtime="00:01:31.12" />
                    <SPLIT distance="200" swimtime="00:02:08.60" />
                    <SPLIT distance="250" swimtime="00:02:37.37" />
                    <SPLIT distance="300" swimtime="00:03:10.11" />
                    <SPLIT distance="350" swimtime="00:03:37.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12408" number="1" />
                    <RELAYPOSITION athleteid="12420" number="2" />
                    <RELAYPOSITION athleteid="12337" number="3" />
                    <RELAYPOSITION athleteid="12371" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="2">
              <RESULTS>
                <RESULT eventid="1122" points="120" swimtime="00:02:45.56" resultid="12459" heatid="12948" lane="2" entrytime="00:02:43.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.30" />
                    <SPLIT distance="100" swimtime="00:01:21.49" />
                    <SPLIT distance="150" swimtime="00:02:05.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12436" number="1" />
                    <RELAYPOSITION athleteid="12384" number="2" />
                    <RELAYPOSITION athleteid="12404" number="3" />
                    <RELAYPOSITION athleteid="12444" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1186" points="354" swimtime="00:04:51.73" resultid="12460" heatid="13041" lane="2" entrytime="00:05:08.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.32" />
                    <SPLIT distance="100" swimtime="00:01:07.15" />
                    <SPLIT distance="150" swimtime="00:01:42.55" />
                    <SPLIT distance="200" swimtime="00:02:24.66" />
                    <SPLIT distance="250" swimtime="00:03:03.03" />
                    <SPLIT distance="300" swimtime="00:03:47.56" />
                    <SPLIT distance="350" swimtime="00:04:17.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12367" number="1" />
                    <RELAYPOSITION athleteid="12428" number="2" />
                    <RELAYPOSITION athleteid="12424" number="3" />
                    <RELAYPOSITION athleteid="12375" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1119" points="133" swimtime="00:03:00.89" resultid="12461" heatid="12946" lane="1" entrytime="00:02:58.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.32" />
                    <SPLIT distance="100" swimtime="00:01:24.43" />
                    <SPLIT distance="150" swimtime="00:02:12.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12341" number="1" />
                    <RELAYPOSITION athleteid="12359" number="2" />
                    <RELAYPOSITION athleteid="12388" number="3" />
                    <RELAYPOSITION athleteid="12363" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SVZ" nation="SUI" region="RZO" clubid="12038" name="Schwimmverein Zürileu" shortname="SV Zürileu">
          <ATHLETES>
            <ATHLETE firstname="Ulises" lastname="Kubli" birthdate="2006-09-12" gender="M" nation="SUI" license="108874" athleteid="13784">
              <RESULTS>
                <RESULT eventid="1141" points="314" swimtime="00:01:11.10" resultid="13785" heatid="12975" lane="1" entrytime="00:01:14.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="298" swimtime="00:01:22.79" resultid="13786" heatid="13017" lane="4" entrytime="00:01:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="David" lastname="Saminskij" birthdate="2007-06-30" gender="M" nation="SUI" license="109445" athleteid="13791">
              <RESULTS>
                <RESULT eventid="1141" points="356" swimtime="00:01:08.14" resultid="13792" heatid="12976" lane="3" entrytime="00:01:12.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="303 - Nicht mit beiden Händen gleichzeitig angeschlagen (Wende  ...)" eventid="1171" status="DSQ" swimtime="00:01:18.22" resultid="13793" heatid="13017" lane="3" entrytime="00:01:20.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Abdurahman" lastname="Serhir" birthdate="2006-05-08" gender="M" nation="SUI" license="20086" athleteid="13794">
              <RESULTS>
                <RESULT eventid="1131" points="275" swimtime="00:01:13.45" resultid="13795" heatid="12959" lane="1" entrytime="00:01:20.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="308" swimtime="00:01:12.96" resultid="13796" heatid="12996" lane="3" entrytime="00:01:12.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Linus" lastname="Bundi" birthdate="2006-09-12" gender="M" nation="SUI" license="122971" athleteid="13781">
              <RESULTS>
                <RESULT eventid="1141" points="276" swimtime="00:01:14.18" resultid="13782" heatid="12975" lane="3" entrytime="00:01:14.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="278" swimtime="00:01:24.78" resultid="13783" heatid="13016" lane="3" entrytime="00:01:27.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dario" lastname="Bundi" birthdate="2006-09-12" gender="M" nation="SUI" license="122972" athleteid="13777">
              <RESULTS>
                <RESULT eventid="1141" points="223" swimtime="00:01:19.58" resultid="13778" heatid="12973" lane="2" entrytime="00:01:22.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="233" swimtime="00:01:29.93" resultid="13779" heatid="13016" lane="4" entrytime="00:01:29.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="306" swimtime="00:01:06.67" resultid="13780" heatid="13037" lane="2" entrytime="00:01:06.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophie" lastname="Kunath" birthdate="2007-08-03" gender="F" nation="SUI" license="108876" athleteid="13787">
              <RESULTS>
                <RESULT eventid="1136" points="343" swimtime="00:01:18.40" resultid="13788" heatid="12966" lane="3" entrytime="00:01:20.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1166" points="364" swimtime="00:01:27.30" resultid="13789" heatid="13011" lane="2" entrytime="00:01:26.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="352" swimtime="00:01:11.16" resultid="13790" heatid="13023" lane="2" entrytime="00:01:11.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1191" points="404" swimtime="00:04:07.42" resultid="13797" heatid="13045" lane="1" entrytime="00:04:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.16" />
                    <SPLIT distance="100" swimtime="00:01:01.09" />
                    <SPLIT distance="150" swimtime="00:01:31.74" />
                    <SPLIT distance="200" swimtime="00:02:04.18" />
                    <SPLIT distance="250" swimtime="00:02:33.94" />
                    <SPLIT distance="300" swimtime="00:03:06.40" />
                    <SPLIT distance="350" swimtime="00:03:35.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13794" number="1" />
                    <RELAYPOSITION athleteid="13784" number="2" />
                    <RELAYPOSITION athleteid="13781" number="3" />
                    <RELAYPOSITION athleteid="13791" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="ALL" nation="SUI" region="RZW" clubid="11839" name="Schwimmclub Allschwil">
          <ATHLETES>
            <ATHLETE firstname="Fabien" lastname="Vogt" birthdate="2001-06-25" gender="M" nation="SUI" license="6395" athleteid="13244">
              <RESULTS>
                <RESULT eventid="1141" points="440" swimtime="00:01:03.50" resultid="13245" heatid="12977" lane="2" entrytime="00:01:01.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="423" swimtime="00:01:05.63" resultid="13246" heatid="12997" lane="3" entrytime="00:01:06.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="468" swimtime="00:00:57.88" resultid="13247" heatid="14655" lane="3" entrytime="00:00:57.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elena" lastname="Geiger" birthdate="2010-03-06" gender="F" nation="SUI" license="32344" athleteid="13221">
              <RESULTS>
                <RESULT comment="304 - Schwimmen in Bauchlage vor der Wende (Wende ...)" eventid="1065" status="DSQ" swimtime="00:01:54.36" resultid="13222" heatid="12857" lane="3" entrytime="00:01:55.40" />
                <RESULT eventid="1099" points="151" swimtime="00:01:56.93" resultid="13223" heatid="12897" lane="3" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="124" swimtime="00:01:40.60" resultid="13224" heatid="12927" lane="2" entrytime="00:01:40.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milo" lastname="Jackson" birthdate="2009-12-11" gender="M" nation="FRA" license="32286" athleteid="13225">
              <RESULTS>
                <RESULT eventid="1070" points="131" swimtime="00:01:35.00" resultid="13226" heatid="12866" lane="2" entrytime="00:01:40.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="160" swimtime="00:01:22.73" resultid="13227" heatid="12939" lane="1" entrytime="00:01:32.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dario" lastname="Meyer" birthdate="2010-07-06" gender="M" nation="SUI" license="6389" athleteid="13232">
              <RESULTS>
                <RESULT eventid="1070" points="87" swimtime="00:01:48.92" resultid="13233" heatid="12865" lane="3" entrytime="00:01:55.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="131" swimtime="00:01:48.85" resultid="13234" heatid="12908" lane="1" entrytime="00:01:57.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="140" swimtime="00:01:26.52" resultid="13235" heatid="12940" lane="1" entrytime="00:01:29.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Lazarevski" birthdate="1999-10-28" gender="M" nation="SUI" license="6404" athleteid="13228">
              <RESULTS>
                <RESULT eventid="1131" points="339" swimtime="00:01:08.51" resultid="13229" heatid="12959" lane="3" entrytime="00:01:17.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="365" swimtime="00:01:08.95" resultid="13230" heatid="12997" lane="4" entrytime="00:01:09.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="389" swimtime="00:01:01.54" resultid="13231" heatid="13040" lane="2" entrytime="00:01:00.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Raphael" lastname="Meyer" birthdate="2012-01-18" gender="M" nation="SUI" license="6429" athleteid="13236">
              <RESULTS>
                <RESULT eventid="1076" points="112" swimtime="00:00:46.07" resultid="13237" heatid="12882" lane="3" entrytime="00:00:48.72" />
                <RESULT eventid="1096" points="99" swimtime="00:00:54.45" resultid="13238" heatid="12894" lane="2" entrytime="00:00:56.88" />
                <RESULT eventid="1109" points="111" swimtime="00:00:41.91" resultid="13239" heatid="12922" lane="1" entrytime="00:00:45.71" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kiara" lastname="Stäheli" birthdate="2010-02-21" gender="F" nation="SUI" license="6410" athleteid="13240">
              <RESULTS>
                <RESULT eventid="1065" points="201" swimtime="00:01:33.65" resultid="13241" heatid="12861" lane="4" entrytime="00:01:41.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="193" swimtime="00:01:26.91" resultid="13242" heatid="12932" lane="1" entrytime="00:01:22.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="162" swimtime="00:01:54.35" resultid="13243" heatid="12901" lane="3" entrytime="00:01:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Camila" lastname="Brugger" birthdate="1999-12-26" gender="F" nation="SUI" license="6384" athleteid="13209">
              <RESULTS>
                <RESULT eventid="1146" points="338" swimtime="00:01:21.06" resultid="13210" heatid="12982" lane="1" entrytime="00:01:26.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="384" swimtime="00:01:09.11" resultid="13211" heatid="13027" lane="1" entrytime="00:01:07.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alvaro" lastname="Cancela" birthdate="2009-02-21" gender="M" nation="SUI" license="6375" athleteid="13212">
              <RESULTS>
                <RESULT eventid="1060" points="200" swimtime="00:00:37.17" resultid="13213" heatid="12854" lane="3" entrytime="00:00:44.78" />
                <RESULT eventid="1070" points="130" swimtime="00:01:35.25" resultid="13214" heatid="12867" lane="3" entrytime="00:01:38.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="183" swimtime="00:01:19.12" resultid="13215" heatid="12940" lane="2" entrytime="00:01:26.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1088" points="175" swimtime="00:02:57.61" resultid="13216" heatid="12884" lane="3" entrytime="00:03:03.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.90" />
                    <SPLIT distance="100" swimtime="00:01:25.53" />
                    <SPLIT distance="150" swimtime="00:02:12.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emilio" lastname="Cancela" birthdate="2012-04-06" gender="M" nation="SUI" license="32276" athleteid="13217">
              <RESULTS>
                <RESULT eventid="1076" points="39" swimtime="00:01:05.26" resultid="13218" heatid="12881" lane="4" entrytime="00:00:59.39" />
                <RESULT eventid="1096" points="62" swimtime="00:01:03.60" resultid="13219" heatid="12894" lane="1" entrytime="00:00:57.46" />
                <RESULT eventid="1109" points="51" swimtime="00:00:54.22" resultid="13220" heatid="12921" lane="3" entrytime="00:00:49.71" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT comment="205 - Frühablösung (Staffelschwimmer ...)" eventid="1122" status="DSQ" swimtime="00:02:33.86" resultid="13248" heatid="14668" lane="1" entrytime="00:02:35.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.27" />
                    <SPLIT distance="100" swimtime="00:01:13.30" />
                    <SPLIT distance="150" swimtime="00:01:58.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13212" number="1" />
                    <RELAYPOSITION athleteid="13232" number="2" />
                    <RELAYPOSITION athleteid="13236" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="13225" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
          <COACHES>
            <COACH firstname="Anja" gender="F" lastname="Bornhauser" license="6380" type="HEADCOACH" />
          </COACHES>
          <OFFICIALS>
            <OFFICIAL officialid="14677" firstname="Brigitte" gender="F" grade="Schiedsrichter" lastname="Feuerbacher" nation="SUI" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="AARE" nation="SUI" region="RZW" clubid="12172" name="Schwimmclub Aarefisch Aarau" shortname="Schwimmclub Aarefisch">
          <ATHLETES>
            <ATHLETE firstname="Sanae" lastname="König" birthdate="2007-07-27" gender="F" nation="SUI" license="110626" athleteid="13130" />
            <ATHLETE firstname="Mailin" lastname="Hösli" birthdate="2007-07-24" gender="F" nation="SUI" license="114230" athleteid="13116">
              <RESULTS>
                <RESULT eventid="1125" points="228" swimtime="00:01:29.31" resultid="13117" heatid="12949" lane="4" entrytime="00:01:39.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="252" swimtime="00:01:26.88" resultid="13118" heatid="12965" lane="1" entrytime="00:01:28.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="259" swimtime="00:01:28.57" resultid="13119" heatid="12980" lane="3" entrytime="00:01:33.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1166" points="274" swimtime="00:01:35.93" resultid="13120" heatid="13010" lane="1" entrytime="00:01:34.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="270" swimtime="00:01:17.67" resultid="13121" heatid="13023" lane="4" entrytime="00:01:13.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yahya" lastname="Hussain" birthdate="2011-03-28" gender="M" nation="SUI" license="123814" athleteid="13122">
              <RESULTS>
                <RESULT eventid="1076" points="92" swimtime="00:00:49.05" resultid="13123" heatid="12879" lane="3" entrytime="00:01:04.99" />
                <RESULT eventid="1096" points="73" swimtime="00:01:00.37" resultid="13124" heatid="12894" lane="4" entrytime="00:01:00.00" />
                <RESULT eventid="1109" points="101" swimtime="00:00:43.25" resultid="13125" heatid="12921" lane="4" entrytime="00:00:52.38" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Luongo" birthdate="2013-05-29" gender="F" nation="SUI" athleteid="13131">
              <RESULTS>
                <RESULT eventid="1073" points="120" swimtime="00:00:51.89" resultid="13132" heatid="12874" lane="1" entrytime="00:00:55.07" />
                <RESULT eventid="1092" points="97" swimtime="00:01:02.01" resultid="13133" heatid="12889" lane="2" entrytime="00:00:59.98" />
                <RESULT eventid="1106" points="141" swimtime="00:00:43.98" resultid="13134" heatid="12916" lane="3" entrytime="00:00:46.82" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giulia" lastname="Morini" birthdate="2006-07-10" gender="F" nation="SUI" license="105646" athleteid="13141">
              <RESULTS>
                <RESULT eventid="1125" points="288" swimtime="00:01:22.61" resultid="13142" heatid="12951" lane="3" entrytime="00:01:24.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="328" swimtime="00:01:19.55" resultid="13143" heatid="12966" lane="2" entrytime="00:01:20.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="310" swimtime="00:01:23.43" resultid="13144" heatid="12984" lane="4" entrytime="00:01:23.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1166" points="211" swimtime="00:01:44.67" resultid="13145" heatid="13009" lane="3" entrytime="00:01:42.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="388" swimtime="00:01:08.86" resultid="13146" heatid="13026" lane="4" entrytime="00:01:08.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="David" lastname="Radam" birthdate="2004-06-06" gender="M" nation="SUI" license="38824" athleteid="13163">
              <RESULTS>
                <RESULT eventid="1131" points="543" swimtime="00:00:58.56" resultid="13164" heatid="14653" lane="2" entrytime="00:00:59.00" />
                <RESULT eventid="1161" points="631" swimtime="00:01:55.82" resultid="13165" heatid="13006" lane="2" entrytime="00:01:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.64" />
                    <SPLIT distance="100" swimtime="00:00:55.86" />
                    <SPLIT distance="150" swimtime="00:01:25.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="551" swimtime="00:00:54.79" resultid="13166" heatid="14655" lane="2" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tobias" lastname="Dietiker" birthdate="2011-09-13" gender="M" nation="SUI" license="123649" athleteid="13092">
              <RESULTS>
                <RESULT eventid="1076" points="92" swimtime="00:00:49.12" resultid="13093" heatid="12882" lane="4" entrytime="00:00:53.87" />
                <RESULT eventid="1096" points="106" swimtime="00:00:53.20" resultid="13094" heatid="12895" lane="1" entrytime="00:00:53.40" />
                <RESULT eventid="1109" points="99" swimtime="00:00:43.48" resultid="13095" heatid="12922" lane="3" entrytime="00:00:43.83" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maksim" lastname="Bucher" birthdate="2013-04-16" gender="M" nation="SUI" license="123651" athleteid="13077">
              <RESULTS>
                <RESULT eventid="1076" points="75" swimtime="00:00:52.49" resultid="13078" heatid="12881" lane="2" entrytime="00:00:54.92" />
                <RESULT eventid="1096" points="59" swimtime="00:01:04.60" resultid="13079" heatid="12892" lane="3" entrytime="00:01:09.61" />
                <RESULT eventid="1109" points="90" swimtime="00:00:44.92" resultid="13080" heatid="12922" lane="4" entrytime="00:00:47.89" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Moira" lastname="Gämperle" birthdate="2011-01-21" gender="F" nation="SUI" athleteid="13101">
              <RESULTS>
                <RESULT eventid="1073" points="156" swimtime="00:00:47.46" resultid="13102" heatid="12877" lane="3" entrytime="00:00:49.35" />
                <RESULT eventid="1092" points="120" swimtime="00:00:57.81" resultid="13103" heatid="12890" lane="4" entrytime="00:00:59.41" />
                <RESULT eventid="1106" points="188" swimtime="00:00:40.02" resultid="13104" heatid="12918" lane="3" entrytime="00:00:41.54" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joshua" lastname="Thölking" birthdate="2009-09-04" gender="M" nation="SUI" license="106821" athleteid="13193">
              <RESULTS>
                <RESULT eventid="1060" points="226" swimtime="00:00:35.70" resultid="13194" heatid="12855" lane="2" entrytime="00:00:37.29" entrycourse="LCM" />
                <RESULT eventid="1070" points="232" swimtime="00:01:18.55" resultid="13195" heatid="12868" lane="2" entrytime="00:01:23.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="222" swimtime="00:01:31.27" resultid="13196" heatid="12910" lane="3" entrytime="00:01:38.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="281" swimtime="00:01:08.60" resultid="13197" heatid="12942" lane="3" entrytime="00:01:11.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lielle" lastname="Jakob" birthdate="2011-06-27" gender="F" nation="SUI" license="121254" athleteid="13126">
              <RESULTS>
                <RESULT eventid="1073" points="108" swimtime="00:00:53.67" resultid="13127" heatid="12874" lane="4" entrytime="00:00:55.07" />
                <RESULT eventid="1092" points="132" swimtime="00:00:56.07" resultid="13128" heatid="12889" lane="3" entrytime="00:00:59.98" />
                <RESULT eventid="1106" points="118" swimtime="00:00:46.67" resultid="13129" heatid="12916" lane="2" entrytime="00:00:46.82" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Soyala" lastname="Deverin" birthdate="2007-10-01" gender="F" nation="SUI" license="121367" athleteid="13086">
              <RESULTS>
                <RESULT eventid="1125" points="334" swimtime="00:01:18.65" resultid="13087" heatid="12952" lane="3" entrytime="00:01:19.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="371" swimtime="00:01:16.33" resultid="13088" heatid="12967" lane="4" entrytime="00:01:18.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="380" swimtime="00:01:17.97" resultid="13089" heatid="12986" lane="1" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1166" points="327" swimtime="00:01:30.44" resultid="13090" heatid="13010" lane="2" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="412" swimtime="00:01:07.50" resultid="13091" heatid="13027" lane="4" entrytime="00:01:07.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Meta" lastname="Zimmermann" birthdate="2006-11-12" gender="F" nation="SUI" license="105340" athleteid="13198">
              <RESULTS>
                <RESULT eventid="1146" points="427" swimtime="00:01:15.02" resultid="13199" heatid="12989" lane="1" entrytime="00:01:14.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="471" swimtime="00:02:21.84" resultid="13200" heatid="13001" lane="4" entrytime="00:02:21.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.09" />
                    <SPLIT distance="100" swimtime="00:01:07.45" />
                    <SPLIT distance="150" swimtime="00:01:44.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="475" swimtime="00:01:04.37" resultid="13201" heatid="13031" lane="4" entrytime="00:01:03.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michelle" lastname="Saxer" birthdate="2007-02-17" gender="F" nation="SUI" license="101862" athleteid="13183">
              <RESULTS>
                <RESULT eventid="1125" points="350" swimtime="00:01:17.43" resultid="13184" heatid="12954" lane="1" entrytime="00:01:15.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="333" swimtime="00:01:19.12" resultid="13185" heatid="12967" lane="1" entrytime="00:01:18.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="318" swimtime="00:01:22.76" resultid="13186" heatid="12987" lane="4" entrytime="00:01:18.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="342" swimtime="00:01:11.80" resultid="13187" heatid="13025" lane="1" entrytime="00:01:09.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alexander" lastname="Hofmann" birthdate="2007-02-14" gender="M" nation="SUI" license="112326" athleteid="13110">
              <RESULTS>
                <RESULT eventid="1131" points="172" swimtime="00:01:25.77" resultid="13111" heatid="12957" lane="1" entrytime="00:01:42.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="169" swimtime="00:01:27.32" resultid="13112" heatid="12970" lane="3" entrytime="00:01:46.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="220" swimtime="00:01:21.61" resultid="13113" heatid="12991" lane="1" entrytime="00:01:38.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="209" swimtime="00:01:33.19" resultid="13114" heatid="13015" lane="1" entrytime="00:01:35.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="290" swimtime="00:01:07.87" resultid="13115" heatid="13038" lane="1" entrytime="00:01:05.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anouk" lastname="Blattner" birthdate="2011-02-16" gender="F" nation="SUI" license="121256" athleteid="13061">
              <RESULTS>
                <RESULT eventid="1073" points="70" swimtime="00:01:01.98" resultid="13062" heatid="12872" lane="4" entrytime="00:01:07.35" />
                <RESULT comment="303 - Nicht mit beiden Händen gleichzeitig angeschlagen (Wende  ...)" eventid="1092" status="DSQ" swimtime="00:00:55.58" resultid="13063" heatid="12891" lane="1" entrytime="00:00:58.70" />
                <RESULT eventid="1106" points="54" swimtime="00:01:00.45" resultid="13064" heatid="12913" lane="4" entrytime="00:00:59.47" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amelia" lastname="Balliello" birthdate="2008-10-28" gender="F" nation="GER" license="121408" athleteid="13051">
              <RESULTS>
                <RESULT eventid="1125" points="193" swimtime="00:01:34.47" resultid="13052" heatid="12949" lane="3" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="183" swimtime="00:01:36.59" resultid="13053" heatid="12962" lane="1" entrytime="00:01:45.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="238" swimtime="00:01:31.14" resultid="13054" heatid="12978" lane="1" entrytime="00:01:48.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1166" points="262" swimtime="00:01:37.41" resultid="13055" heatid="13010" lane="4" entrytime="00:01:41.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="214" swimtime="00:01:23.97" resultid="13056" heatid="13019" lane="2" entrytime="00:01:25.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Samantha" lastname="Stucki" birthdate="2010-04-20" gender="F" nation="SUI" athleteid="13188">
              <RESULTS>
                <RESULT eventid="1099" points="144" swimtime="00:01:58.93" resultid="13189" heatid="12897" lane="2" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="231" swimtime="00:01:21.83" resultid="13190" heatid="12928" lane="3" entrytime="00:01:30.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1053" points="153" swimtime="00:00:45.58" resultid="13191" heatid="12847" lane="2" entrytime="00:00:50.25" />
                <RESULT eventid="1065" points="193" swimtime="00:01:34.89" resultid="13192" heatid="12860" lane="2" entrytime="00:01:41.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Michelle" lastname="Armandi" birthdate="2006-11-20" gender="F" nation="SUI" athleteid="13046">
              <RESULTS>
                <RESULT eventid="1125" points="482" swimtime="00:01:09.62" resultid="13047" heatid="12954" lane="3" entrytime="00:01:12.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="487" swimtime="00:01:11.81" resultid="13048" heatid="12987" lane="2" entrytime="00:01:17.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="574" swimtime="00:02:12.83" resultid="13049" heatid="13001" lane="3" entrytime="00:02:18.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.36" />
                    <SPLIT distance="100" swimtime="00:01:05.47" />
                    <SPLIT distance="150" swimtime="00:01:40.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="534" swimtime="00:01:01.92" resultid="13050" heatid="13031" lane="2" entrytime="00:01:02.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Noemi" lastname="Nguyen" birthdate="2008-12-31" gender="F" nation="SUI" license="120934" athleteid="13147">
              <RESULTS>
                <RESULT eventid="1125" status="WDR" swimtime="00:00:00.00" resultid="13148" entrytime="00:01:23.50" entrycourse="LCM" />
                <RESULT eventid="1136" status="WDR" swimtime="00:00:00.00" resultid="13149" entrytime="00:01:27.26" entrycourse="LCM" />
                <RESULT eventid="1146" status="WDR" swimtime="00:00:00.00" resultid="13150" entrytime="00:01:39.42" entrycourse="SCM" />
                <RESULT eventid="1166" status="WDR" swimtime="00:00:00.00" resultid="13151" entrytime="00:01:33.65" entrycourse="LCM" />
                <RESULT eventid="1176" status="WDR" swimtime="00:00:00.00" resultid="13152" entrytime="00:01:13.01" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andreina" lastname="Hoffmann" birthdate="2010-05-24" gender="F" nation="SUI" license="112378" athleteid="13105">
              <RESULTS>
                <RESULT eventid="1053" status="WDR" swimtime="00:00:00.00" resultid="13106" heatid="12849" lane="4" entrytime="00:00:46.93" />
                <RESULT eventid="1065" status="WDR" swimtime="00:00:00.00" resultid="13107" heatid="12862" lane="4" entrytime="00:01:35.05" />
                <RESULT eventid="1099" status="WDR" swimtime="00:00:00.00" resultid="13108" heatid="12899" lane="2" entrytime="00:01:53.88" />
                <RESULT eventid="1112" status="WDR" swimtime="00:00:00.00" resultid="13109" heatid="12932" lane="4" entrytime="00:01:22.21" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yannick" lastname="Rohr" birthdate="2006-12-05" gender="M" nation="SUI" license="114844" athleteid="13173">
              <RESULTS>
                <RESULT eventid="1131" points="255" swimtime="00:01:15.33" resultid="13174" heatid="12959" lane="2" entrytime="00:01:16.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="257" swimtime="00:01:16.01" resultid="13175" heatid="12974" lane="3" entrytime="00:01:20.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="310" swimtime="00:01:12.79" resultid="13176" heatid="12996" lane="4" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="269" swimtime="00:01:25.70" resultid="13177" heatid="13015" lane="2" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="348" swimtime="00:01:03.86" resultid="13178" heatid="13038" lane="3" entrytime="00:01:04.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Noé Alexander" lastname="Bolliger" birthdate="2004-12-08" gender="M" nation="SUI" license="47174" athleteid="13065">
              <RESULTS>
                <RESULT eventid="1131" status="WDR" swimtime="00:00:00.00" resultid="13066" heatid="12960" lane="1" entrytime="00:01:14.67" entrycourse="LCM" />
                <RESULT eventid="1141" status="WDR" swimtime="00:00:00.00" resultid="13067" heatid="12975" lane="4" entrytime="00:01:16.07" entrycourse="SCM" />
                <RESULT eventid="1151" status="WDR" swimtime="00:00:00.00" resultid="13068" heatid="12996" lane="1" entrytime="00:01:14.21" entrycourse="SCM" />
                <RESULT eventid="1171" status="WDR" swimtime="00:00:00.00" resultid="13069" heatid="13017" lane="2" entrytime="00:01:17.12" entrycourse="LCM" />
                <RESULT eventid="1181" status="WDR" swimtime="00:00:00.00" resultid="13070" heatid="13040" lane="3" entrytime="00:01:00.77" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manon" lastname="Bircher" birthdate="2011-04-24" gender="F" nation="SUI" athleteid="13057">
              <RESULTS>
                <RESULT eventid="1073" status="WDR" swimtime="00:00:00.00" resultid="13058" heatid="12877" lane="1" entrytime="00:00:49.73" />
                <RESULT eventid="1092" status="WDR" swimtime="00:00:00.00" resultid="13059" heatid="14113" lane="1" entrytime="00:00:53.83" />
                <RESULT eventid="1106" status="WDR" swimtime="00:00:00.00" resultid="13060" heatid="12918" lane="4" entrytime="00:00:43.19" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabian" lastname="Radam" birthdate="2008-07-06" gender="M" nation="GER" license="109621" athleteid="13167">
              <RESULTS>
                <RESULT eventid="1131" points="237" swimtime="00:01:17.17" resultid="13168" heatid="12958" lane="1" entrytime="00:01:22.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="322" swimtime="00:01:10.49" resultid="13169" heatid="12976" lane="2" entrytime="00:01:12.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="292" swimtime="00:01:14.28" resultid="13170" heatid="12994" lane="4" entrytime="00:01:23.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="268" swimtime="00:01:25.79" resultid="13171" heatid="13016" lane="1" entrytime="00:01:29.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="301" swimtime="00:01:07.04" resultid="13172" heatid="13037" lane="4" entrytime="00:01:08.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Danyal" lastname="Nisamov" birthdate="2010-07-18" gender="M" nation="SUI" license="119001" athleteid="13153">
              <RESULTS>
                <RESULT eventid="1070" points="101" swimtime="00:01:43.69" resultid="13154" heatid="12867" lane="1" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="95" swimtime="00:02:00.87" resultid="13155" heatid="12908" lane="4" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="103" swimtime="00:01:35.63" resultid="13156" heatid="12940" lane="4" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emilie" lastname="Sandberg" birthdate="2011-05-16" gender="F" nation="SWE" license="120921" athleteid="13179">
              <RESULTS>
                <RESULT eventid="1073" points="116" swimtime="00:00:52.43" resultid="13180" heatid="12873" lane="1" entrytime="00:00:57.93" />
                <RESULT comment="303 - Nicht mit beiden Händen gleichzeitig angeschlagen (Wende  ...)" eventid="1092" status="DSQ" swimtime="00:01:01.91" resultid="13181" heatid="12887" lane="3" entrytime="00:01:06.23" />
                <RESULT eventid="1106" points="149" swimtime="00:00:43.16" resultid="13182" heatid="12917" lane="2" entrytime="00:00:43.84" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emeline" lastname="Durrieu" birthdate="2011-05-25" gender="F" nation="SUI" athleteid="13096">
              <RESULTS>
                <RESULT eventid="1073" points="85" swimtime="00:00:58.02" resultid="13097" heatid="12873" lane="3" entrytime="00:00:57.89" />
                <RESULT eventid="1092" points="121" swimtime="00:00:57.68" resultid="13098" heatid="12888" lane="2" entrytime="00:01:00.33" />
                <RESULT eventid="1106" points="118" swimtime="00:00:46.62" resultid="13099" heatid="12917" lane="3" entrytime="00:00:44.73" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lars" lastname="Oeschger" birthdate="2007-09-11" gender="M" nation="SUI" license="106711" athleteid="13157">
              <RESULTS>
                <RESULT eventid="1131" points="264" swimtime="00:01:14.42" resultid="13158" heatid="12960" lane="3" entrytime="00:01:14.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="232" swimtime="00:01:18.55" resultid="13159" heatid="12973" lane="3" entrytime="00:01:22.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="255" swimtime="00:01:17.63" resultid="13160" heatid="12992" lane="2" entrytime="00:01:27.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="223" swimtime="00:01:31.24" resultid="13161" heatid="13013" lane="2" entrytime="00:01:44.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="291" swimtime="00:01:07.81" resultid="13162" heatid="13037" lane="3" entrytime="00:01:07.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Flavia" lastname="Gjata" birthdate="2008-12-22" gender="F" nation="SUI" license="122582" athleteid="13100">
              <RESULTS>
                <RESULT eventid="1125" status="WDR" swimtime="00:00:00.00" resultid="14050" heatid="12950" lane="1" entrytime="00:01:30.00" />
                <RESULT eventid="1166" status="WDR" swimtime="00:00:00.00" resultid="14051" heatid="13009" lane="1" entrytime="00:01:44.64" />
                <RESULT eventid="1146" status="WDR" swimtime="00:00:00.00" resultid="14052" heatid="12980" lane="1" entrytime="00:01:35.00" />
                <RESULT eventid="1176" status="WDR" swimtime="00:00:00.00" resultid="14054" heatid="13022" lane="2" entrytime="00:01:14.75" />
                <RESULT eventid="1136" status="WDR" swimtime="00:00:00.00" resultid="14055" heatid="12964" lane="3" entrytime="00:01:31.88" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dario" lastname="Boxler" birthdate="2005-05-24" gender="M" nation="SUI" license="38808" athleteid="13071">
              <RESULTS>
                <RESULT eventid="1131" points="382" swimtime="00:01:05.81" resultid="13072" heatid="14653" lane="4" entrytime="00:01:09.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="354" swimtime="00:01:08.32" resultid="13073" heatid="12976" lane="4" entrytime="00:01:12.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="403" swimtime="00:01:06.68" resultid="13074" heatid="12996" lane="2" entrytime="00:01:09.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="443" swimtime="00:01:12.57" resultid="13075" heatid="13018" lane="2" entrytime="00:01:11.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="382" swimtime="00:01:01.93" resultid="13076" heatid="14655" lane="4" entrytime="00:00:59.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hanna" lastname="Meier" birthdate="2008-07-06" gender="F" nation="SUI" license="114409" athleteid="13135">
              <RESULTS>
                <RESULT eventid="1125" points="157" swimtime="00:01:41.04" resultid="13136" heatid="12949" lane="1" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="246" swimtime="00:01:27.55" resultid="13137" heatid="12964" lane="2" entrytime="00:01:31.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="264" swimtime="00:01:28.02" resultid="13138" heatid="12979" lane="1" entrytime="00:01:39.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1166" points="261" swimtime="00:01:37.56" resultid="13139" heatid="13009" lane="2" entrytime="00:01:41.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="281" swimtime="00:01:16.71" resultid="13140" heatid="13022" lane="1" entrytime="00:01:16.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stella" lastname="Campbell" birthdate="2010-10-24" gender="F" nation="SUI" license="121275" athleteid="13081">
              <RESULTS>
                <RESULT eventid="1053" points="160" swimtime="00:00:44.90" resultid="13082" heatid="12848" lane="2" entrytime="00:00:47.96" />
                <RESULT eventid="1065" points="218" swimtime="00:01:31.18" resultid="13083" heatid="12862" lane="3" entrytime="00:01:34.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="171" swimtime="00:01:52.29" resultid="13084" heatid="12902" lane="3" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="221" swimtime="00:01:22.99" resultid="13085" heatid="12929" lane="3" entrytime="00:01:27.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1122" points="137" swimtime="00:02:38.50" resultid="13202" heatid="12948" lane="3" entrytime="00:02:49.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.09" />
                    <SPLIT distance="100" swimtime="00:01:23.10" />
                    <SPLIT distance="150" swimtime="00:02:06.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13153" number="1" />
                    <RELAYPOSITION athleteid="13122" number="2" />
                    <RELAYPOSITION athleteid="13092" number="3" />
                    <RELAYPOSITION athleteid="13193" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1191" points="411" swimtime="00:04:06.07" resultid="13203" heatid="13045" lane="3" entrytime="00:04:04.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.72" />
                    <SPLIT distance="100" swimtime="00:01:05.08" />
                    <SPLIT distance="150" swimtime="00:01:36.55" />
                    <SPLIT distance="200" swimtime="00:02:12.16" />
                    <SPLIT distance="250" swimtime="00:02:40.49" />
                    <SPLIT distance="300" swimtime="00:03:11.51" />
                    <SPLIT distance="350" swimtime="00:03:37.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13173" number="1" />
                    <RELAYPOSITION athleteid="13110" number="2" />
                    <RELAYPOSITION athleteid="13071" number="3" />
                    <RELAYPOSITION athleteid="13163" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1119" points="194" swimtime="00:02:39.52" resultid="13204" heatid="12946" lane="2" entrytime="00:02:31.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.38" />
                    <SPLIT distance="100" swimtime="00:01:18.11" />
                    <SPLIT distance="150" swimtime="00:01:54.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13188" number="1" />
                    <RELAYPOSITION athleteid="13101" number="2" />
                    <RELAYPOSITION athleteid="13081" number="3" />
                    <RELAYPOSITION athleteid="13096" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1186" points="437" swimtime="00:04:31.96" resultid="13205" heatid="13042" lane="3" entrytime="00:04:39.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.34" />
                    <SPLIT distance="100" swimtime="00:01:07.09" />
                    <SPLIT distance="150" swimtime="00:01:39.71" />
                    <SPLIT distance="200" swimtime="00:02:16.29" />
                    <SPLIT distance="250" swimtime="00:02:47.34" />
                    <SPLIT distance="300" swimtime="00:03:21.67" />
                    <SPLIT distance="350" swimtime="00:03:55.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13086" number="1" />
                    <RELAYPOSITION athleteid="13141" number="2" />
                    <RELAYPOSITION athleteid="13198" number="3" />
                    <RELAYPOSITION athleteid="13183" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1119" points="115" swimtime="00:03:10.02" resultid="13206" heatid="12945" lane="2" entrytime="00:03:15.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.69" />
                    <SPLIT distance="100" swimtime="00:01:42.94" />
                    <SPLIT distance="150" swimtime="00:02:26.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13179" number="1" />
                    <RELAYPOSITION athleteid="13061" number="2" />
                    <RELAYPOSITION athleteid="13131" number="3" />
                    <RELAYPOSITION athleteid="13126" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1186" points="315" swimtime="00:05:03.42" resultid="13207" heatid="13042" lane="1" entrytime="00:04:56.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.41" />
                    <SPLIT distance="100" swimtime="00:01:01.92" />
                    <SPLIT distance="150" swimtime="00:01:37.38" />
                    <SPLIT distance="200" swimtime="00:02:19.22" />
                    <SPLIT distance="250" swimtime="00:02:55.88" />
                    <SPLIT distance="300" swimtime="00:03:37.43" />
                    <SPLIT distance="350" swimtime="00:04:16.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13046" number="1" />
                    <RELAYPOSITION athleteid="13135" number="2" />
                    <RELAYPOSITION athleteid="13116" number="3" />
                    <RELAYPOSITION athleteid="13051" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
          <COACHES>
            <COACH firstname="Piotr" gender="M" lastname="Albinski" nation="POL" type="HEADCOACH" />
          </COACHES>
        </CLUB>
        <CLUB type="CLUB" code="REG" nation="SUI" region="RZO" clubid="12782" name="Schwimmclub Regensdorf" shortname="Scr">
          <ATHLETES>
            <ATHLETE firstname="Moira" lastname="Steiner" birthdate="2007-08-10" gender="F" nation="SUI" license="113684" athleteid="14157">
              <RESULTS>
                <RESULT comment="209 - Zehen beider Füsse nicht in Kontakt mit Wand oder Anschlagplatte (Start)" eventid="1136" status="DSQ" swimtime="00:01:21.12" resultid="14158" heatid="12967" lane="2" entrytime="00:01:18.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1166" points="295" swimtime="00:01:33.59" resultid="14159" heatid="13011" lane="4" entrytime="00:01:29.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="374" swimtime="00:01:09.72" resultid="14160" heatid="13028" lane="3" entrytime="00:01:06.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="318" swimtime="00:01:22.74" resultid="14161" heatid="12981" lane="4" entrytime="00:01:30.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="324" swimtime="00:02:40.69" resultid="14162" heatid="12998" lane="1" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.32" />
                    <SPLIT distance="100" swimtime="00:01:16.90" />
                    <SPLIT distance="150" swimtime="00:01:59.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kilian" lastname="Dell&apos; Agosti" birthdate="2012-10-04" gender="M" nation="SUI" athleteid="14121">
              <RESULTS>
                <RESULT eventid="1076" points="63" swimtime="00:00:55.75" resultid="14122" heatid="12880" lane="1" entrytime="00:01:01.21" entrycourse="SCM" />
                <RESULT eventid="1096" points="75" swimtime="00:00:59.64" resultid="14123" heatid="12893" lane="3" entrytime="00:01:03.93" entrycourse="SCM" />
                <RESULT eventid="1109" points="60" swimtime="00:00:51.23" resultid="14124" heatid="12920" lane="1" entrytime="00:00:56.72" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nora" lastname="Zurbuchen" birthdate="2009-08-22" gender="F" nation="SUI" athleteid="14163">
              <RESULTS>
                <RESULT eventid="1065" points="177" swimtime="00:01:37.62" resultid="14164" heatid="12860" lane="1" entrytime="00:01:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="254" swimtime="00:01:38.34" resultid="14165" heatid="12899" lane="4" entrytime="00:01:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="176" swimtime="00:01:29.53" resultid="14166" heatid="12929" lane="1" entrytime="00:01:28.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natasha" lastname="Kaluperuma de Silva" birthdate="2009-01-31" gender="F" nation="SUI" athleteid="14146">
              <RESULTS>
                <RESULT eventid="1084" points="242" swimtime="00:02:57.11" resultid="14147" heatid="12883" lane="2" entrytime="00:03:00.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.05" />
                    <SPLIT distance="100" swimtime="00:01:28.07" />
                    <SPLIT distance="150" swimtime="00:02:13.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="247" swimtime="00:01:20.03" resultid="14148" heatid="12932" lane="3" entrytime="00:01:21.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Selina" lastname="Dürler" birthdate="2011-06-27" gender="F" nation="SUI" athleteid="14138">
              <RESULTS>
                <RESULT eventid="1073" points="189" swimtime="00:00:44.55" resultid="14139" heatid="12877" lane="2" entrytime="00:00:48.58" entrycourse="SCM" />
                <RESULT eventid="1092" points="151" swimtime="00:00:53.59" resultid="14140" heatid="14113" lane="4" entrytime="00:00:55.47" entrycourse="SCM" />
                <RESULT eventid="1106" points="179" swimtime="00:00:40.68" resultid="14141" heatid="12918" lane="1" entrytime="00:00:41.88" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kevin" lastname="Dell&apos; Agosti" birthdate="2009-09-13" gender="M" nation="SUI" license="124393" athleteid="14116">
              <RESULTS>
                <RESULT eventid="1060" points="74" swimtime="00:00:51.72" resultid="14117" heatid="12853" lane="4" entrytime="00:00:54.48" entrycourse="SCM" />
                <RESULT eventid="1070" points="98" swimtime="00:01:44.63" resultid="14118" heatid="12866" lane="1" entrytime="00:01:43.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="133" swimtime="00:01:48.29" resultid="14119" heatid="12908" lane="2" entrytime="00:01:53.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="107" swimtime="00:01:34.39" resultid="14120" heatid="12939" lane="4" entrytime="00:01:33.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kirsten" lastname="Roso" birthdate="2008-06-26" gender="F" nation="INA" license="117429" athleteid="14153">
              <RESULTS>
                <RESULT eventid="1146" points="204" swimtime="00:01:35.85" resultid="14154" heatid="12979" lane="2" entrytime="00:01:35.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="191" swimtime="00:01:27.17" resultid="14155" heatid="13020" lane="3" entrytime="00:01:23.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1166" points="191" swimtime="00:01:48.23" resultid="14156" heatid="13008" lane="2" entrytime="00:01:45.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marianna" lastname="Dohmen" birthdate="2009-03-20" gender="F" nation="SUI" license="121732" athleteid="14129">
              <RESULTS>
                <RESULT eventid="1099" points="200" swimtime="00:01:46.57" resultid="14130" heatid="12900" lane="2" entrytime="00:01:52.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1065" points="168" swimtime="00:01:39.45" resultid="14131" heatid="12856" lane="3" />
                <RESULT eventid="1112" points="136" swimtime="00:01:37.53" resultid="14132" heatid="12925" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Christina" lastname="Dohmen" birthdate="2010-11-03" gender="F" nation="SUI" license="121731" athleteid="14125">
              <RESULTS>
                <RESULT eventid="1065" points="127" swimtime="00:01:49.10" resultid="14126" heatid="12858" lane="2" entrytime="00:01:51.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="148" swimtime="00:01:57.82" resultid="14127" heatid="12898" lane="2" entrytime="00:01:57.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="125" swimtime="00:01:40.42" resultid="14128" heatid="12927" lane="3" entrytime="00:01:41.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vincent Luis" lastname="Küppers" birthdate="2013-01-29" gender="M" nation="GER" athleteid="14149">
              <RESULTS>
                <RESULT comment="304 - Schwimmen in Bauchlage vor der Wende (Wende ...)" eventid="1076" status="DSQ" swimtime="00:00:59.20" resultid="14150" heatid="12880" lane="3" entrytime="00:01:00.97" entrycourse="SCM" />
                <RESULT comment="525 - Füsse während der Vortriebsphase nicht nach aussen gedreht" eventid="1096" status="DSQ" swimtime="00:01:06.30" resultid="14151" heatid="12892" lane="2" entrytime="00:01:06.72" entrycourse="SCM" />
                <RESULT eventid="1109" points="68" swimtime="00:00:49.16" resultid="14152" heatid="12921" lane="2" entrytime="00:00:49.54" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Niklas" lastname="Grabenweger" birthdate="2011-10-02" gender="M" nation="AUT" athleteid="14142">
              <RESULTS>
                <RESULT eventid="1076" points="52" swimtime="00:00:59.42" resultid="14143" heatid="12879" lane="2" entrytime="00:01:04.11" entrycourse="SCM" />
                <RESULT eventid="1096" points="67" swimtime="00:01:01.94" resultid="14144" heatid="12893" lane="4" entrytime="00:01:06.34" entrycourse="SCM" />
                <RESULT eventid="1109" points="75" swimtime="00:00:47.69" resultid="14145" heatid="12920" lane="2" entrytime="00:00:53.06" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amanda" lastname="Dürler" birthdate="2008-07-06" gender="F" nation="SUI" license="120217" athleteid="14133">
              <RESULTS>
                <RESULT eventid="1136" points="225" swimtime="00:01:30.15" resultid="14134" heatid="12965" lane="4" entrytime="00:01:29.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="203" swimtime="00:01:36.15" resultid="14135" heatid="12978" lane="3" entrytime="00:01:41.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1166" points="158" swimtime="00:01:55.17" resultid="14136" heatid="13007" lane="1" entrytime="00:01:52.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="236" swimtime="00:01:21.20" resultid="14137" heatid="13022" lane="4" entrytime="00:01:17.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1122" points="78" swimtime="00:03:10.91" resultid="14665" heatid="12947" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.26" />
                    <SPLIT distance="100" swimtime="00:01:39.93" />
                    <SPLIT distance="150" swimtime="00:02:29.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14116" number="1" />
                    <RELAYPOSITION athleteid="14121" number="2" />
                    <RELAYPOSITION athleteid="14142" number="3" />
                    <RELAYPOSITION athleteid="14149" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1119" points="196" swimtime="00:02:38.98" resultid="14666" heatid="12944" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.83" />
                    <SPLIT distance="100" swimtime="00:01:25.88" />
                    <SPLIT distance="150" swimtime="00:02:02.72" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="14146" number="1" />
                    <RELAYPOSITION athleteid="14125" number="2" />
                    <RELAYPOSITION athleteid="14138" number="3" />
                    <RELAYPOSITION athleteid="14163" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="BIRS" nation="SUI" region="RZW" clubid="12816" name="Schwimmclub Birsfelden" shortname="Scbirs">
          <ATHLETES>
            <ATHLETE firstname="Cilia" lastname="Jeker" birthdate="2008-03-20" gender="F" nation="SUI" athleteid="13417">
              <RESULTS>
                <RESULT eventid="1136" points="211" swimtime="00:01:32.15" resultid="13418" heatid="12964" lane="4" entrytime="00:01:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="237" swimtime="00:01:31.29" resultid="13419" heatid="12981" lane="3" entrytime="00:01:29.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="245" swimtime="00:01:20.21" resultid="13420" heatid="13021" lane="4" entrytime="00:01:19.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alina" lastname="Sturzenegger" birthdate="2008-06-26" gender="F" nation="SUI" athleteid="13432">
              <RESULTS>
                <RESULT eventid="1136" points="230" swimtime="00:01:29.58" resultid="13433" heatid="12964" lane="1" entrytime="00:01:34.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="251" swimtime="00:01:29.54" resultid="13434" heatid="12982" lane="4" entrytime="00:01:27.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="264" swimtime="00:01:18.27" resultid="13435" heatid="13021" lane="3" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jan" lastname="Stalder" birthdate="2010-06-28" gender="M" nation="SUI" athleteid="13430">
              <RESULTS>
                <RESULT eventid="1116" status="WDR" swimtime="00:00:00.00" resultid="13431" heatid="12936" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alexandra Nina" lastname="van Dongen" birthdate="2006-05-20" gender="F" nation="SUI" athleteid="13439">
              <RESULTS>
                <RESULT eventid="1136" points="125" swimtime="00:01:49.77" resultid="13440" heatid="12962" lane="2" entrytime="00:01:44.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="164" swimtime="00:01:31.71" resultid="13441" heatid="13020" lane="4" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksa" lastname="Zivanovic" birthdate="2010-12-21" gender="M" nation="SUI" athleteid="13442">
              <RESULTS>
                <RESULT eventid="1070" points="94" swimtime="00:01:45.92" resultid="13443" heatid="12864" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="82" swimtime="00:01:43.31" resultid="13444" heatid="12936" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Naomi" lastname="Klopfstein" birthdate="2004-08-17" gender="F" nation="SUI" athleteid="13421">
              <RESULTS>
                <RESULT comment="306 - Wand in Bauchlage verlassen  (Wende ...)" eventid="1136" status="DSQ" swimtime="00:01:59.92" resultid="13422" heatid="12963" lane="1" entrytime="00:01:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="164" swimtime="00:01:31.74" resultid="13423" heatid="13020" lane="1" entrytime="00:01:24.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valentin" lastname="Tschopp" birthdate="2010-04-07" gender="M" nation="SUI" athleteid="13436">
              <RESULTS>
                <RESULT eventid="1070" points="33" swimtime="00:02:29.38" resultid="13437" heatid="12864" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="43" swimtime="00:02:07.66" resultid="13438" heatid="12936" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Morris" lastname="Reetz" birthdate="2008-06-30" gender="M" nation="SUI" athleteid="13427">
              <RESULTS>
                <RESULT eventid="1141" points="80" swimtime="00:01:52.12" resultid="13428" heatid="12971" lane="1" entrytime="00:01:43.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="110" swimtime="00:01:33.52" resultid="13429" heatid="13033" lane="3" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pascual" lastname="Mencìa" birthdate="2010-12-18" gender="F" nation="SUI" athleteid="13424">
              <RESULTS>
                <RESULT comment="404 - Nicht in Rückenlage angeschlagen (Ziel)" eventid="1065" status="DSQ" swimtime="00:01:51.73" resultid="13425" heatid="12856" lane="1" />
                <RESULT eventid="1112" points="171" swimtime="00:01:30.47" resultid="13426" heatid="12925" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1186" points="216" swimtime="00:05:44.10" resultid="13445" heatid="13041" lane="3" entrytime="00:05:23.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.10" />
                    <SPLIT distance="100" swimtime="00:01:22.63" />
                    <SPLIT distance="150" swimtime="00:02:04.16" />
                    <SPLIT distance="200" swimtime="00:02:54.55" />
                    <SPLIT distance="250" swimtime="00:03:37.46" />
                    <SPLIT distance="300" swimtime="00:04:25.58" />
                    <SPLIT distance="350" swimtime="00:05:02.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13417" number="1" />
                    <RELAYPOSITION athleteid="13421" number="2" />
                    <RELAYPOSITION athleteid="13439" number="3" />
                    <RELAYPOSITION athleteid="13432" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="LIES" nation="SUI" region="RZW" clubid="12060" name="Schwimmclub Liestal">
          <ATHLETES>
            <ATHLETE firstname="Céline" lastname="Müller" birthdate="2006-08-17" gender="F" nation="SUI" license="104766" athleteid="13515">
              <RESULTS>
                <RESULT eventid="1136" points="502" swimtime="00:01:09.03" resultid="13516" heatid="12969" lane="3" entrytime="00:01:09.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="369" swimtime="00:01:18.75" resultid="13517" heatid="12989" lane="4" entrytime="00:01:15.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fiona Valentina" lastname="Flückiger" birthdate="2010-04-09" gender="F" nation="SUI" license="115257" athleteid="13476">
              <RESULTS>
                <RESULT eventid="1053" points="239" swimtime="00:00:39.25" resultid="13477" heatid="12850" lane="2" entrytime="00:00:40.31" entrycourse="LCM" />
                <RESULT eventid="1099" points="243" swimtime="00:01:39.82" resultid="13478" heatid="12902" lane="2" entrytime="00:01:44.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="242" swimtime="00:01:20.55" resultid="13479" heatid="12930" lane="1" entrytime="00:01:25.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alexander" lastname="Wacker" birthdate="2010-05-25" gender="M" nation="GER" athleteid="13545">
              <RESULTS>
                <RESULT eventid="1103" points="97" swimtime="00:02:00.38" resultid="13546" heatid="12906" lane="2" entrytime="00:02:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="39" swimtime="00:02:11.57" resultid="13547" heatid="12937" lane="3" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lia" lastname="Schiess" birthdate="2006-08-25" gender="F" nation="SUI" license="7933" athleteid="13539">
              <RESULTS>
                <RESULT eventid="1136" points="455" swimtime="00:01:11.35" resultid="13540" heatid="12969" lane="4" entrytime="00:01:11.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="493" swimtime="00:01:03.58" resultid="13541" heatid="13031" lane="3" entrytime="00:01:03.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lena" lastname="Gessesse" birthdate="2010-03-09" gender="F" nation="SUI" license="119428" athleteid="13480">
              <RESULTS>
                <RESULT eventid="1053" points="235" swimtime="00:00:39.49" resultid="13481" heatid="12850" lane="3" entrytime="00:00:40.72" entrycourse="LCM" />
                <RESULT eventid="1065" points="230" swimtime="00:01:29.57" resultid="13482" heatid="12862" lane="1" entrytime="00:01:34.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="227" swimtime="00:01:22.29" resultid="13483" heatid="12930" lane="3" entrytime="00:01:24.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Xenia" lastname="Blumin" birthdate="2006-09-30" gender="F" nation="SUI" license="115281" athleteid="13462">
              <RESULTS>
                <RESULT eventid="1146" points="520" swimtime="00:01:10.24" resultid="13463" heatid="12990" lane="2" entrytime="00:01:09.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1166" points="426" swimtime="00:01:22.82" resultid="13464" heatid="13012" lane="2" entrytime="00:01:22.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="598" swimtime="00:01:05.14" resultid="14672" heatid="12969" lane="2" entrytime="00:01:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lennon" lastname="Schmied" birthdate="2007-08-17" gender="M" nation="SUI" license="111478" athleteid="13542">
              <RESULTS>
                <RESULT eventid="1141" points="216" swimtime="00:01:20.47" resultid="13543" heatid="12973" lane="1" entrytime="00:01:25.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1161" points="265" swimtime="00:02:34.66" resultid="13544" heatid="13004" lane="3" entrytime="00:02:38.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.88" />
                    <SPLIT distance="100" swimtime="00:01:17.11" />
                    <SPLIT distance="150" swimtime="00:01:58.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giordana" lastname="Graf" birthdate="2008-08-20" gender="F" nation="SUI" license="105829" athleteid="13484">
              <RESULTS>
                <RESULT eventid="1125" points="317" swimtime="00:01:20.03" resultid="13485" heatid="12951" lane="2" entrytime="00:01:23.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="398" swimtime="00:01:16.77" resultid="13486" heatid="12981" lane="2" entrytime="00:01:28.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1166" points="415" swimtime="00:01:23.60" resultid="13487" heatid="13012" lane="4" entrytime="00:01:25.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Max" lastname="Saxer" birthdate="2009-09-10" gender="M" nation="SUI" athleteid="13532">
              <RESULTS>
                <RESULT comment="206 - Unterwasserphase: Mehr als ein Delphinbeinschlag (Start)" eventid="1103" status="DSQ" swimtime="00:01:59.63" resultid="13533" heatid="12906" lane="3" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="41" swimtime="00:02:09.44" resultid="13534" heatid="12937" lane="2" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rebekka" lastname="Jäger" birthdate="2009-08-02" gender="F" nation="SUI" license="111475" athleteid="13491">
              <RESULTS>
                <RESULT eventid="1053" points="236" swimtime="00:00:39.43" resultid="13492" heatid="12849" lane="3" entrytime="00:00:42.29" entrycourse="LCM" />
                <RESULT eventid="1084" points="349" swimtime="00:02:36.80" resultid="13493" heatid="14112" lane="1" entrytime="00:02:48.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.70" />
                    <SPLIT distance="100" swimtime="00:01:14.55" />
                    <SPLIT distance="150" swimtime="00:01:55.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="360" swimtime="00:01:10.58" resultid="13494" heatid="12934" lane="2" entrytime="00:01:11.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julie Pascale" lastname="Räuber" birthdate="2009-03-18" gender="F" nation="SUI" license="119430" athleteid="13525">
              <RESULTS>
                <RESULT eventid="1065" points="219" swimtime="00:01:30.93" resultid="13526" heatid="12863" lane="4" entrytime="00:01:27.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.37" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="204 - Starten vor dem Startkommando" eventid="1099" status="DSQ" swimtime="00:01:41.26" resultid="13527" heatid="12903" lane="4" entrytime="00:01:42.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="270" swimtime="00:01:17.74" resultid="13528" heatid="12933" lane="3" entrytime="00:01:16.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fiona" lastname="Liesch" birthdate="2006-06-07" gender="F" nation="SUI" license="100547" athleteid="13505">
              <RESULTS>
                <RESULT eventid="1156" points="527" swimtime="00:02:16.67" resultid="13506" heatid="13001" lane="1" entrytime="00:02:20.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.07" />
                    <SPLIT distance="100" swimtime="00:01:05.12" />
                    <SPLIT distance="150" swimtime="00:01:40.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="474" swimtime="00:01:12.43" resultid="13507" heatid="12990" lane="4" entrytime="00:01:12.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1166" points="492" swimtime="00:01:18.97" resultid="14671" heatid="14115" lane="2" entrytime="00:01:16.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kilian" lastname="Roppel" birthdate="2007-02-09" gender="M" nation="SUI" license="100566" athleteid="13529">
              <RESULTS>
                <RESULT eventid="1151" points="236" swimtime="00:01:19.67" resultid="13530" heatid="12993" lane="4" entrytime="00:01:25.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="221" swimtime="00:01:14.32" resultid="13531" heatid="13038" lane="4" entrytime="00:01:06.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Melanie" lastname="Allemann" birthdate="2010-01-01" gender="F" nation="SUI" license="111473" athleteid="13446">
              <RESULTS>
                <RESULT comment="302 - Wand nicht berührt (Wende ...)" eventid="1065" status="DSQ" swimtime="00:01:34.65" resultid="13447" heatid="12861" lane="3" entrytime="00:01:38.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="244" swimtime="00:01:39.67" resultid="13448" heatid="12902" lane="1" entrytime="00:01:45.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="215" swimtime="00:01:23.79" resultid="13449" heatid="12930" lane="4" entrytime="00:01:25.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Severin" lastname="Oberli" birthdate="2007-09-28" gender="M" nation="SUI" license="104767" athleteid="13522">
              <RESULTS>
                <RESULT eventid="1141" points="298" swimtime="00:01:12.34" resultid="13523" heatid="12974" lane="2" entrytime="00:01:17.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1161" points="300" swimtime="00:02:28.31" resultid="13524" heatid="13005" lane="1" entrytime="00:02:32.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.34" />
                    <SPLIT distance="100" swimtime="00:01:11.26" />
                    <SPLIT distance="150" swimtime="00:01:50.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolas" lastname="Nietschmann" birthdate="2006-08-30" gender="M" nation="SUI" license="115623" athleteid="13518">
              <RESULTS>
                <RESULT eventid="1131" points="387" swimtime="00:01:05.52" resultid="13519" heatid="14653" lane="3" entrytime="00:01:04.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="345" swimtime="00:01:10.21" resultid="13520" heatid="12995" lane="2" entrytime="00:01:15.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="368" swimtime="00:01:02.71" resultid="13521" heatid="13039" lane="4" entrytime="00:01:03.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yannick" lastname="Knab" birthdate="2006-05-09" gender="M" nation="SUI" license="100563" athleteid="13498">
              <RESULTS>
                <RESULT eventid="1141" points="355" swimtime="00:01:08.20" resultid="13499" heatid="12976" lane="1" entrytime="00:01:12.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1161" points="366" swimtime="00:02:18.81" resultid="13500" heatid="13005" lane="2" entrytime="00:02:25.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.29" />
                    <SPLIT distance="100" swimtime="00:01:06.26" />
                    <SPLIT distance="150" swimtime="00:01:43.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ellie" lastname="Wartenweiler" birthdate="2008-07-04" gender="F" nation="SUI" license="123105" athleteid="13548">
              <RESULTS>
                <RESULT eventid="1146" points="301" swimtime="00:01:24.28" resultid="13549" heatid="12980" lane="4" entrytime="00:01:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1166" points="218" swimtime="00:01:43.57" resultid="13550" heatid="13007" lane="3" entrytime="00:01:52.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="298" swimtime="00:01:15.18" resultid="13551" heatid="13021" lane="2" entrytime="00:01:17.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Talia" lastname="Jordan" birthdate="2007-06-06" gender="F" nation="SUI" license="105237" athleteid="13495">
              <RESULTS>
                <RESULT eventid="1146" points="516" swimtime="00:01:10.44" resultid="13496" heatid="12988" lane="3" entrytime="00:01:16.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="506" swimtime="00:01:03.05" resultid="13497" heatid="13031" lane="1" entrytime="00:01:03.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Layra" lastname="Balmer" birthdate="2009-03-15" gender="F" nation="SUI" license="115255" athleteid="13450">
              <RESULTS>
                <RESULT eventid="1053" points="303" swimtime="00:00:36.28" resultid="13451" heatid="12851" lane="1" entrytime="00:00:39.75" entrycourse="LCM" />
                <RESULT eventid="1084" points="337" swimtime="00:02:38.57" resultid="13452" heatid="14112" lane="2" entrytime="00:02:44.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.02" />
                    <SPLIT distance="100" swimtime="00:01:15.27" />
                    <SPLIT distance="150" swimtime="00:01:57.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="359" swimtime="00:01:10.65" resultid="13453" heatid="12934" lane="1" entrytime="00:01:13.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Camille" lastname="Schicktanz" birthdate="2009-07-05" gender="F" nation="SUI" license="111477" athleteid="13535">
              <RESULTS>
                <RESULT eventid="1053" points="325" swimtime="00:00:35.46" resultid="13536" heatid="12851" lane="2" entrytime="00:00:36.04" entrycourse="LCM" />
                <RESULT eventid="1084" points="303" swimtime="00:02:44.26" resultid="13537" heatid="14112" lane="3" entrytime="00:02:47.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.79" />
                    <SPLIT distance="100" swimtime="00:01:19.61" />
                    <SPLIT distance="150" swimtime="00:02:03.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="317" swimtime="00:01:13.69" resultid="13538" heatid="12934" lane="4" entrytime="00:01:15.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Hinnerks" birthdate="2004-12-27" gender="F" nation="SUI" license="117024" athleteid="13488">
              <RESULTS>
                <RESULT eventid="1146" points="483" swimtime="00:01:12.01" resultid="13489" heatid="12990" lane="3" entrytime="00:01:09.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1166" points="474" swimtime="00:01:19.94" resultid="13490" heatid="14115" lane="3" entrytime="00:01:18.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anine" lastname="Ecoffey" birthdate="2010-10-21" gender="F" nation="SUI" license="112809" athleteid="13469">
              <RESULTS>
                <RESULT eventid="1053" points="211" swimtime="00:00:40.92" resultid="13470" heatid="12850" lane="4" entrytime="00:00:41.24" entrycourse="LCM" />
                <RESULT eventid="1099" points="298" swimtime="00:01:33.36" resultid="13471" heatid="12904" lane="4" entrytime="00:01:38.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="256" swimtime="00:01:19.08" resultid="13472" heatid="12933" lane="4" entrytime="00:01:20.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sarina" lastname="Liesch" birthdate="2003-08-09" gender="F" nation="SUI" license="36137" athleteid="13508">
              <RESULTS>
                <RESULT eventid="1136" status="WDR" swimtime="00:00:00.00" resultid="13509" entrytime="00:01:10.62" entrycourse="SCM" />
                <RESULT eventid="1166" status="WDR" swimtime="00:00:00.00" resultid="13510" entrytime="00:01:14.25" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Léna" lastname="Ecoffey" birthdate="2007-12-24" gender="F" nation="SUI" license="105228" athleteid="13473">
              <RESULTS>
                <RESULT eventid="1125" points="520" swimtime="00:01:07.87" resultid="13474" heatid="12955" lane="3" entrytime="00:01:09.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="536" swimtime="00:01:09.56" resultid="13475" heatid="12988" lane="4" entrytime="00:01:17.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dascha" lastname="Blumin" birthdate="2009-02-22" gender="F" nation="SUI" license="123827" athleteid="13458">
              <RESULTS>
                <RESULT eventid="1065" points="300" swimtime="00:01:21.92" resultid="13459" heatid="12863" lane="1" entrytime="00:01:24.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="277" swimtime="00:01:35.57" resultid="13460" heatid="12903" lane="3" entrytime="00:01:39.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="297" swimtime="00:01:15.30" resultid="13461" heatid="12933" lane="1" entrytime="00:01:18.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Flavia" lastname="Meier" birthdate="2008-08-31" gender="F" nation="SUI" license="115259" athleteid="13511">
              <RESULTS>
                <RESULT eventid="1146" points="266" swimtime="00:01:27.81" resultid="13512" heatid="12979" lane="4" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1166" points="238" swimtime="00:01:40.62" resultid="13513" heatid="13008" lane="1" entrytime="00:01:45.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="267" swimtime="00:01:17.96" resultid="13514" heatid="13021" lane="1" entrytime="00:01:18.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna-Maxie" lastname="Leupin" birthdate="2011-05-15" gender="F" nation="SUI" athleteid="13501">
              <RESULTS>
                <RESULT eventid="1073" points="116" swimtime="00:00:52.49" resultid="13502" heatid="12873" lane="4" entrytime="00:00:58.00" />
                <RESULT eventid="1092" points="133" swimtime="00:00:55.95" resultid="13503" heatid="12890" lane="3" entrytime="00:00:59.00" />
                <RESULT eventid="1106" points="136" swimtime="00:00:44.58" resultid="13504" heatid="12914" lane="4" entrytime="00:00:52.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ryan" lastname="Balmer" birthdate="2010-05-18" gender="M" nation="SUI" license="115256" athleteid="13454">
              <RESULTS>
                <RESULT eventid="1070" points="161" swimtime="00:01:28.75" resultid="13455" heatid="12868" lane="1" entrytime="00:01:27.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="141" swimtime="00:01:46.10" resultid="13456" heatid="12910" lane="4" entrytime="00:01:49.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="183" swimtime="00:01:19.09" resultid="13457" heatid="12941" lane="2" entrytime="00:01:18.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" number="1">
              <RESULTS>
                <RESULT eventid="1191" points="328" swimtime="00:04:25.22" resultid="13552" heatid="13044" lane="3" entrytime="00:04:26.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.79" />
                    <SPLIT distance="100" swimtime="00:01:02.29" />
                    <SPLIT distance="150" swimtime="00:01:36.16" />
                    <SPLIT distance="200" swimtime="00:02:13.44" />
                    <SPLIT distance="250" swimtime="00:02:45.37" />
                    <SPLIT distance="300" swimtime="00:03:21.29" />
                    <SPLIT distance="350" swimtime="00:03:51.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13518" number="1" />
                    <RELAYPOSITION athleteid="13542" number="2" />
                    <RELAYPOSITION athleteid="13522" number="3" />
                    <RELAYPOSITION athleteid="13498" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1119" points="366" swimtime="00:02:09.24" resultid="13553" heatid="14669" lane="2" entrytime="00:02:10.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                    <SPLIT distance="100" swimtime="00:01:04.79" />
                    <SPLIT distance="150" swimtime="00:01:36.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13491" number="1" />
                    <RELAYPOSITION athleteid="13450" number="2" />
                    <RELAYPOSITION athleteid="13535" number="3" />
                    <RELAYPOSITION athleteid="13525" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" number="1">
              <RESULTS>
                <RESULT eventid="1186" points="562" swimtime="00:04:10.20" resultid="13554" heatid="13043" lane="2" entrytime="00:04:07.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.58" />
                    <SPLIT distance="100" swimtime="00:01:02.62" />
                    <SPLIT distance="150" swimtime="00:01:32.09" />
                    <SPLIT distance="200" swimtime="00:02:05.39" />
                    <SPLIT distance="250" swimtime="00:02:35.57" />
                    <SPLIT distance="300" swimtime="00:03:08.51" />
                    <SPLIT distance="350" swimtime="00:03:37.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13462" number="1" />
                    <RELAYPOSITION athleteid="13488" number="2" />
                    <RELAYPOSITION athleteid="13505" number="3" />
                    <RELAYPOSITION athleteid="13473" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1119" points="273" swimtime="00:02:22.51" resultid="13555" heatid="14669" lane="1" entrytime="00:02:23.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.93" />
                    <SPLIT distance="100" swimtime="00:01:09.32" />
                    <SPLIT distance="150" swimtime="00:01:46.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13458" number="1" />
                    <RELAYPOSITION athleteid="13469" number="2" />
                    <RELAYPOSITION athleteid="13476" number="3" />
                    <RELAYPOSITION athleteid="13480" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" number="2">
              <RESULTS>
                <RESULT eventid="1186" points="519" swimtime="00:04:16.99" resultid="13556" heatid="13043" lane="1" entrytime="00:04:12.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.42" />
                    <SPLIT distance="100" swimtime="00:01:04.88" />
                    <SPLIT distance="150" swimtime="00:01:35.96" />
                    <SPLIT distance="200" swimtime="00:02:08.65" />
                    <SPLIT distance="250" swimtime="00:02:38.66" />
                    <SPLIT distance="300" swimtime="00:03:11.71" />
                    <SPLIT distance="350" swimtime="00:03:43.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="13539" number="1" />
                    <RELAYPOSITION athleteid="13515" number="2" />
                    <RELAYPOSITION athleteid="13495" number="3" />
                    <RELAYPOSITION athleteid="13484" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SCUW" nation="SUI" region="RZO" clubid="12462" name="Schwimmclub Uster Wallisellen" shortname="SC Uster Wallisellen">
          <ATHLETES>
            <ATHLETE firstname="Samuele" lastname="Di Toffa" birthdate="2006-12-26" gender="M" nation="SUI" license="103620" athleteid="13607">
              <RESULTS>
                <RESULT eventid="1131" points="287" swimtime="00:01:12.36" resultid="13608" heatid="12960" lane="4" entrytime="00:01:15.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="295" swimtime="00:01:14.01" resultid="13609" heatid="12994" lane="2" entrytime="00:01:18.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="382" swimtime="00:01:01.89" resultid="13610" heatid="13038" lane="2" entrytime="00:01:03.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Krista" lastname="Fischer" birthdate="2003-08-24" gender="F" nation="GER" license="100584" athleteid="13611">
              <RESULTS>
                <RESULT eventid="1136" points="346" swimtime="00:01:18.17" resultid="13612" heatid="12968" lane="1" entrytime="00:01:14.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="358" swimtime="00:01:19.53" resultid="13613" heatid="12987" lane="1" entrytime="00:01:18.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1166" points="320" swimtime="00:01:31.09" resultid="13614" heatid="13011" lane="1" entrytime="00:01:29.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valentina" lastname="Nocito" birthdate="2005-03-22" gender="F" nation="SUI" license="107794" athleteid="13615">
              <RESULTS>
                <RESULT eventid="1125" status="SICK" swimtime="00:00:00.00" resultid="13616" heatid="12952" lane="1" entrytime="00:01:19.83" entrycourse="SCM" />
                <RESULT eventid="1146" status="SICK" swimtime="00:00:00.00" resultid="13617" heatid="12985" lane="2" entrytime="00:01:20.68" entrycourse="SCM" />
                <RESULT eventid="1176" status="SICK" swimtime="00:00:00.00" resultid="13618" heatid="13025" lane="2" entrytime="00:01:09.16" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Moritz" lastname="Kessler" birthdate="2003-12-26" gender="M" nation="SUI" athleteid="14167">
              <RESULTS>
                <RESULT eventid="1151" points="251" swimtime="00:01:18.10" resultid="14168" heatid="12995" lane="1" entrytime="00:01:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="266" swimtime="00:01:26.03" resultid="14169" heatid="13016" lane="2" entrytime="00:01:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1181" points="305" swimtime="00:01:06.69" resultid="14170" heatid="13036" lane="3" entrytime="00:01:11.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sinja" lastname="Steinegger" birthdate="2005-10-11" gender="F" nation="SUI" license="103930" athleteid="13619">
              <RESULTS>
                <RESULT eventid="1136" status="WDR" swimtime="00:00:00.00" resultid="13620" heatid="12968" lane="3" entrytime="00:01:12.94" entrycourse="LCM" />
                <RESULT eventid="1146" status="WDR" swimtime="00:00:00.00" resultid="13621" heatid="12988" lane="2" entrytime="00:01:16.26" entrycourse="SCM" />
                <RESULT eventid="1166" status="WDR" swimtime="00:00:00.00" resultid="13622" heatid="13012" lane="1" entrytime="00:01:25.46" entrycourse="SCM" />
                <RESULT eventid="1176" status="WDR" swimtime="00:00:00.00" resultid="13623" heatid="13029" lane="3" entrytime="00:01:05.03" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
  <TIMESTANDARDLISTS>
    <TIMESTANDARDLIST timestandardlistid="5605" course="SCM" gender="M" name="Fricktalcup 2013 Nachmittag" type="MAXIMUM">
      <AGEGROUP agemax="-1" agemin="13" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:35.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="5607" course="SCM" gender="F" name="Fricktalcup 2013 Nachmittag" type="MAXIMUM">
      <AGEGROUP agemax="-1" agemin="13" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:35.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="5601" course="SCM" gender="M" name="Fricktalcup 2013 Vormittag" type="MAXIMUM">
      <AGEGROUP agemax="12" agemin="-1" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:00:55.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:17.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="5603" course="SCM" gender="F" name="Fricktalcup 2013 Vormittag" type="MAXIMUM">
      <AGEGROUP agemax="12" agemin="-1" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:00:55.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:17.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
  </TIMESTANDARDLISTS>
</LENEX>
